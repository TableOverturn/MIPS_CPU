/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : vga_sec_ram                                                  **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module vga_sec_ram( CLK,
                    LOGISIM_CLOCK_TREE_0,
                    R0,
                    R1,
                    R2,
                    R3,
                    R4,
                    R5,
                    R6,
                    R7,
                    R8,
                    R9,
                    R10,
                    R11,
                    R12,
                    R13,
                    R14,
                    R15,
                    Write,
                    input_X,
                    addr,
                    bit_out);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input  CLK;
   input[4:0]  LOGISIM_CLOCK_TREE_0;
   input[31:0]  R0;
   input[31:0]  R1;
   input[31:0]  R2;
   input[31:0]  R3;
   input[31:0]  R4;
   input[31:0]  R5;
   input[31:0]  R6;
   input[31:0]  R7;
   input[31:0]  R8;
   input[31:0]  R9;
   input[31:0]  R10;
   input[31:0]  R11;
   input[31:0]  R12;
   input[31:0]  R13;
   input[31:0]  R14;
   input[31:0]  R15;

   input  Write;
   input[3:0]  input_X;
   input[8:0]  addr;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output bit_out;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   wire[3:0] s_LOGISIM_BUS_10;
   wire[3:0] s_LOGISIM_BUS_101;
   wire[31:0] s_LOGISIM_BUS_102;
   wire[3:0] s_LOGISIM_BUS_104;
   wire[3:0] s_LOGISIM_BUS_107;
   wire[3:0] s_LOGISIM_BUS_108;
   wire[3:0] s_LOGISIM_BUS_109;
   wire[31:0] s_LOGISIM_BUS_11;
   wire[3:0] s_LOGISIM_BUS_110;
   wire[3:0] s_LOGISIM_BUS_111;
   wire[3:0] s_LOGISIM_BUS_113;
   wire[3:0] s_LOGISIM_BUS_114;
   wire[3:0] s_LOGISIM_BUS_115;
   wire[3:0] s_LOGISIM_BUS_116;
   wire[3:0] s_LOGISIM_BUS_119;
   wire[3:0] s_LOGISIM_BUS_120;
   wire[3:0] s_LOGISIM_BUS_21;
   wire[31:0] s_LOGISIM_BUS_24;
   wire[3:0] s_LOGISIM_BUS_27;
   wire[31:0] s_LOGISIM_BUS_30;
   wire[8:0] s_LOGISIM_BUS_35;
   wire[31:0] s_LOGISIM_BUS_39;
   wire[3:0] s_LOGISIM_BUS_40;
   wire[31:0] s_LOGISIM_BUS_49;
   wire[31:0] s_LOGISIM_BUS_5;
   wire[3:0] s_LOGISIM_BUS_50;
   wire[31:0] s_LOGISIM_BUS_51;
   wire[31:0] s_LOGISIM_BUS_53;
   wire[31:0] s_LOGISIM_BUS_57;
   wire[31:0] s_LOGISIM_BUS_58;
   wire[31:0] s_LOGISIM_BUS_6;
   wire[3:0] s_LOGISIM_BUS_60;
   wire[31:0] s_LOGISIM_BUS_67;
   wire[3:0] s_LOGISIM_BUS_68;
   wire[3:0] s_LOGISIM_BUS_70;
   wire[3:0] s_LOGISIM_BUS_72;
   wire[3:0] s_LOGISIM_BUS_74;
   wire[3:0] s_LOGISIM_BUS_75;
   wire[31:0] s_LOGISIM_BUS_8;
   wire[31:0] s_LOGISIM_BUS_82;
   wire[3:0] s_LOGISIM_BUS_83;
   wire[3:0] s_LOGISIM_BUS_85;
   wire[3:0] s_LOGISIM_BUS_88;
   wire[3:0] s_LOGISIM_BUS_89;
   wire[3:0] s_LOGISIM_BUS_90;
   wire[3:0] s_LOGISIM_BUS_92;
   wire[3:0] s_LOGISIM_BUS_93;
   wire[3:0] s_LOGISIM_BUS_96;
   wire[31:0] s_LOGISIM_BUS_97;
   wire[31:0] s_LOGISIM_BUS_98;
   wire[3:0] s_LOGISIM_BUS_99;
   wire s_LOGISIM_NET_0;
   wire s_LOGISIM_NET_100;
   wire s_LOGISIM_NET_105;
   wire s_LOGISIM_NET_112;
   wire s_LOGISIM_NET_118;
   wire s_LOGISIM_NET_121;
   wire s_LOGISIM_NET_122;
   wire s_LOGISIM_NET_14;
   wire s_LOGISIM_NET_16;
   wire s_LOGISIM_NET_17;
   wire s_LOGISIM_NET_22;
   wire s_LOGISIM_NET_25;
   wire s_LOGISIM_NET_26;
   wire s_LOGISIM_NET_28;
   wire s_LOGISIM_NET_29;
   wire s_LOGISIM_NET_3;
   wire s_LOGISIM_NET_32;
   wire s_LOGISIM_NET_34;
   wire s_LOGISIM_NET_37;
   wire s_LOGISIM_NET_42;
   wire s_LOGISIM_NET_43;
   wire s_LOGISIM_NET_47;
   wire s_LOGISIM_NET_54;
   wire s_LOGISIM_NET_56;
   wire s_LOGISIM_NET_61;
   wire s_LOGISIM_NET_62;
   wire s_LOGISIM_NET_63;
   wire s_LOGISIM_NET_64;
   wire s_LOGISIM_NET_69;
   wire s_LOGISIM_NET_7;
   wire s_LOGISIM_NET_76;
   wire s_LOGISIM_NET_77;
   wire s_LOGISIM_NET_78;
   wire s_LOGISIM_NET_81;
   wire s_LOGISIM_NET_84;
   wire s_LOGISIM_NET_87;
   wire s_LOGISIM_NET_94;
   wire s_LOGISIM_NET_95;


   /***************************************************************************
    ** Here all input connections are defined                                **
    ***************************************************************************/
   assign s_LOGISIM_BUS_97[31:0]             = R5;
   assign s_LOGISIM_BUS_98[31:0]             = R15;
   assign s_LOGISIM_NET_122                  = CLK;
   assign s_LOGISIM_BUS_57[31:0]             = R4;
   assign s_LOGISIM_BUS_39[31:0]             = R1;
   assign s_LOGISIM_BUS_58[31:0]             = R12;
   assign s_LOGISIM_BUS_51[31:0]             = R14;
   assign s_LOGISIM_BUS_24[31:0]             = R7;
   assign s_LOGISIM_BUS_6[31:0]              = R3;
   assign s_LOGISIM_BUS_82[31:0]             = R0;
   assign s_LOGISIM_BUS_53[31:0]             = R9;
   assign s_LOGISIM_BUS_49[31:0]             = R2;
   assign s_LOGISIM_BUS_5[31:0]              = R6;
   assign s_LOGISIM_BUS_11[31:0]             = R13;
   assign s_LOGISIM_BUS_30[31:0]             = R11;
   assign s_LOGISIM_BUS_119[3:0]             = input_X;
   assign s_LOGISIM_NET_121                  = Write;
   assign s_LOGISIM_BUS_67[31:0]             = R10;
   assign s_LOGISIM_BUS_8[31:0]              = R8;
   assign s_LOGISIM_BUS_35[8:0]              = addr;

   /***************************************************************************
    ** Here all output connections are defined                               **
    ***************************************************************************/
   assign bit_out                            = s_LOGISIM_NET_94;

   /***************************************************************************
    ** Here all in-lined components are defined                              **
    ***************************************************************************/
   assign s_LOGISIM_NET_112 = 1'd0;


   /***************************************************************************
    ** Here all normal components are defined                                **
    ***************************************************************************/
   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_1 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
             .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
             .MuxOut(s_LOGISIM_BUS_10[3:0]),
             .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_2 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
             .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
             .MuxOut(s_LOGISIM_BUS_99[3:0]),
             .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_1 (.addr(s_LOGISIM_BUS_115[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[0]),
                                  .q(s_LOGISIM_NET_87),
                                  .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_2 (.addr(s_LOGISIM_BUS_85[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[9]),
                                  .q(s_LOGISIM_NET_17),
                                  .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_3 (.addr(s_LOGISIM_BUS_70[3:0]),
                                 .clk(s_LOGISIM_NET_122),
                                 .d(s_LOGISIM_BUS_102[22]),
                                 .q(s_LOGISIM_NET_16),
                                 .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_4 (.addr(s_LOGISIM_BUS_109[3:0]),
                                 .clk(s_LOGISIM_NET_122),
                                 .d(s_LOGISIM_BUS_102[29]),
                                 .q(s_LOGISIM_NET_61),
                                 .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_3 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
             .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
             .MuxOut(s_LOGISIM_BUS_60[3:0]),
             .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_4 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
             .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
             .MuxOut(s_LOGISIM_BUS_40[3:0]),
             .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_5 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
             .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
             .MuxOut(s_LOGISIM_BUS_120[3:0]),
             .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_6 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
             .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
             .MuxOut(s_LOGISIM_BUS_96[3:0]),
             .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_7 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
             .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
             .MuxOut(s_LOGISIM_BUS_50[3:0]),
             .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_5 (.addr(s_LOGISIM_BUS_111[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[16]),
                                  .q(s_LOGISIM_NET_43),
                                  .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_6 (.addr(s_LOGISIM_BUS_113[3:0]),
                                 .clk(s_LOGISIM_NET_122),
                                 .d(s_LOGISIM_BUS_102[25]),
                                 .q(s_LOGISIM_NET_95),
                                 .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_8 (.Enable(1'b1),
             .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
             .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
             .MuxOut(s_LOGISIM_BUS_68[3:0]),
             .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_7 (.addr(s_LOGISIM_BUS_68[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[15]),
                                  .q(s_LOGISIM_NET_14),
                                  .we(s_LOGISIM_NET_121));

   Multiplexer_2      MUX_9 (.Enable(1'b1),
                             .MuxIn_0(s_LOGISIM_NET_112),
                             .MuxIn_1(s_LOGISIM_NET_100),
                             .MuxOut(s_LOGISIM_NET_94),
                             .Sel(s_LOGISIM_NET_118));

   RAM_vga_sec_ram      RAM_8 (.addr(s_LOGISIM_BUS_83[3:0]),
                                 .clk(s_LOGISIM_NET_122),
                                 .d(s_LOGISIM_BUS_102[27]),
                                 .q(s_LOGISIM_NET_28),
                                 .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_10 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_113[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_11 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_74[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_12 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_85[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_9 (.addr(s_LOGISIM_BUS_116[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[5]),
                                  .q(s_LOGISIM_NET_84),
                                  .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_10 (.addr(s_LOGISIM_BUS_90[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[2]),
                                   .q(s_LOGISIM_NET_64),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_11 (.addr(s_LOGISIM_BUS_40[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[4]),
                                   .q(s_LOGISIM_NET_47),
                                   .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_13 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_21[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_14 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_93[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_15 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_110[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_16 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_83[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_12 (.addr(s_LOGISIM_BUS_75[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[18]),
                                   .q(s_LOGISIM_NET_37),
                                   .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_17 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_90[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_16 #(.NrOfBits(32))
      MUX_18 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_82[31:0]),
              .MuxIn_1(s_LOGISIM_BUS_39[31:0]),
              .MuxIn_10(s_LOGISIM_BUS_67[31:0]),
              .MuxIn_11(s_LOGISIM_BUS_30[31:0]),
              .MuxIn_12(s_LOGISIM_BUS_58[31:0]),
              .MuxIn_13(s_LOGISIM_BUS_11[31:0]),
              .MuxIn_14(s_LOGISIM_BUS_51[31:0]),
              .MuxIn_15(s_LOGISIM_BUS_98[31:0]),
              .MuxIn_2(s_LOGISIM_BUS_49[31:0]),
              .MuxIn_3(s_LOGISIM_BUS_6[31:0]),
              .MuxIn_4(s_LOGISIM_BUS_57[31:0]),
              .MuxIn_5(s_LOGISIM_BUS_97[31:0]),
              .MuxIn_6(s_LOGISIM_BUS_5[31:0]),
              .MuxIn_7(s_LOGISIM_BUS_24[31:0]),
              .MuxIn_8(s_LOGISIM_BUS_8[31:0]),
              .MuxIn_9(s_LOGISIM_BUS_53[31:0]),
              .MuxOut(s_LOGISIM_BUS_102[31:0]),
              .Sel(s_LOGISIM_BUS_119[3:0]));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_19 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_104[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_20 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_107[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_13 (.addr(s_LOGISIM_BUS_114[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[12]),
                                   .q(s_LOGISIM_NET_25),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_14 (.addr(s_LOGISIM_BUS_60[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[10]),
                                   .q(s_LOGISIM_NET_7),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_15 (.addr(s_LOGISIM_BUS_110[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[6]),
                                   .q(s_LOGISIM_NET_54),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_16 (.addr(s_LOGISIM_BUS_101[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[8]),
                                   .q(s_LOGISIM_NET_3),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_17 (.addr(s_LOGISIM_BUS_93[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[30]),
                                  .q(s_LOGISIM_NET_69),
                                  .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_18 (.addr(s_LOGISIM_BUS_89[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[14]),
                                   .q(s_LOGISIM_NET_32),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_19 (.addr(s_LOGISIM_BUS_88[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[21]),
                                   .q(s_LOGISIM_NET_56),
                                   .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_21 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_109[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_22 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_92[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_23 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_101[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_24 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_114[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_25 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_75[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_20 (.addr(s_LOGISIM_BUS_10[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[24]),
                                  .q(s_LOGISIM_NET_34),
                                  .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_21 (.addr(s_LOGISIM_BUS_21[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[11]),
                                   .q(s_LOGISIM_NET_26),
                                   .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_26 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_89[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_27 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_88[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_22 (.addr(s_LOGISIM_BUS_99[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[26]),
                                  .q(s_LOGISIM_NET_78),
                                  .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_28 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_72[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_23 (.addr(s_LOGISIM_BUS_50[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[19]),
                                   .q(s_LOGISIM_NET_63),
                                   .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_29 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_27[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_24 (.addr(s_LOGISIM_BUS_107[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[20]),
                                   .q(s_LOGISIM_NET_77),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_25 (.addr(s_LOGISIM_BUS_96[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[17]),
                                   .q(s_LOGISIM_NET_22),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_26 (.addr(s_LOGISIM_BUS_92[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[7]),
                                   .q(s_LOGISIM_NET_0),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_27 (.addr(s_LOGISIM_BUS_104[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[13]),
                                   .q(s_LOGISIM_NET_62),
                                   .we(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_28 (.addr(s_LOGISIM_BUS_120[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[28]),
                                  .q(s_LOGISIM_NET_81),
                                  .we(s_LOGISIM_NET_121));

   Multiplexer_32      MUX_30 (.Enable(1'b1),
                               .MuxIn_0(s_LOGISIM_NET_29),
                               .MuxIn_1(s_LOGISIM_NET_69),
                               .MuxIn_10(s_LOGISIM_NET_56),
                               .MuxIn_11(s_LOGISIM_NET_77),
                               .MuxIn_12(s_LOGISIM_NET_63),
                               .MuxIn_13(s_LOGISIM_NET_37),
                               .MuxIn_14(s_LOGISIM_NET_22),
                               .MuxIn_15(s_LOGISIM_NET_43),
                               .MuxIn_16(s_LOGISIM_NET_14),
                               .MuxIn_17(s_LOGISIM_NET_32),
                               .MuxIn_18(s_LOGISIM_NET_62),
                               .MuxIn_19(s_LOGISIM_NET_25),
                               .MuxIn_2(s_LOGISIM_NET_61),
                               .MuxIn_20(s_LOGISIM_NET_26),
                               .MuxIn_21(s_LOGISIM_NET_7),
                               .MuxIn_22(s_LOGISIM_NET_17),
                               .MuxIn_23(s_LOGISIM_NET_3),
                               .MuxIn_24(s_LOGISIM_NET_0),
                               .MuxIn_25(s_LOGISIM_NET_54),
                               .MuxIn_26(s_LOGISIM_NET_84),
                               .MuxIn_27(s_LOGISIM_NET_47),
                               .MuxIn_28(s_LOGISIM_NET_105),
                               .MuxIn_29(s_LOGISIM_NET_64),
                               .MuxIn_3(s_LOGISIM_NET_81),
                               .MuxIn_30(s_LOGISIM_NET_42),
                               .MuxIn_31(s_LOGISIM_NET_87),
                               .MuxIn_4(s_LOGISIM_NET_28),
                               .MuxIn_5(s_LOGISIM_NET_78),
                               .MuxIn_6(s_LOGISIM_NET_95),
                               .MuxIn_7(s_LOGISIM_NET_34),
                               .MuxIn_8(s_LOGISIM_NET_76),
                               .MuxIn_9(s_LOGISIM_NET_16),
                               .MuxOut(s_LOGISIM_NET_100),
                               .Sel(s_LOGISIM_BUS_35[8:4]));

   NOT_GATE      GATE_1 (.Input_1(s_LOGISIM_NET_121),
                         .Result(s_LOGISIM_NET_118));

   RAM_vga_sec_ram      RAM_29 (.addr(s_LOGISIM_BUS_74[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[31]),
                                  .q(s_LOGISIM_NET_29),
                                  .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_31 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_115[3:0]),
              .Sel(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_32 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_116[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_30 (.addr(s_LOGISIM_BUS_108[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[1]),
                                   .q(s_LOGISIM_NET_42),
                                   .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_33 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_111[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_31 (.addr(s_LOGISIM_BUS_27[3:0]),
                                  .clk(s_LOGISIM_NET_122),
                                  .d(s_LOGISIM_BUS_102[23]),
                                  .q(s_LOGISIM_NET_76),
                                  .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_34 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_108[3:0]),
              .Sel(s_LOGISIM_NET_121));

   RAM_vga_sec_ram      RAM_32 (.addr(s_LOGISIM_BUS_72[3:0]),
                                   .clk(s_LOGISIM_NET_122),
                                   .d(s_LOGISIM_BUS_102[3]),
                                   .q(s_LOGISIM_NET_105),
                                   .we(s_LOGISIM_NET_121));

   Multiplexer_bus_2 #(.NrOfBits(4))
      MUX_35 (.Enable(1'b1),
              .MuxIn_0(s_LOGISIM_BUS_35[3:0]),
              .MuxIn_1(s_LOGISIM_BUS_119[3:0]),
              .MuxOut(s_LOGISIM_BUS_70[3:0]),
              .Sel(s_LOGISIM_NET_121));



endmodule
