/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : ctrl_sig_autogen                                             **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module ctrl_sig_autogen( F0,
                         F1,
                         F2,
                         F3,
                         F4,
                         F5,
                         LOGISIM_CLOCK_TREE_0,
                         OP0,
                         OP1,
                         OP2,
                         OP3,
                         OP4,
                         OP5,
                         ALU_SRC,
                         BEQ,
                         BLEZ,
                         BNE,
                         HalfW,
                         JAL,
                         JR,
                         JUMP,
                         MemToReg,
                         MemWrite,
                         RegDst,
                         RegWrite,
                         SignedExt,
                         SysCALL,
                         Vshamt);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input  F0;
   input  F1;
   input  F2;
   input  F3;
   input  F4;
   input  F5;
   input[4:0]  LOGISIM_CLOCK_TREE_0;
   input  OP0;
   input  OP1;
   input  OP2;
   input  OP3;
   input  OP4;
   input  OP5;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output ALU_SRC;
   output BEQ;
   output BLEZ;
   output BNE;
   output HalfW;
   output JAL;
   output JR;
   output JUMP;
   output MemToReg;
   output MemWrite;
   output RegDst;
   output RegWrite;
   output SignedExt;
   output SysCALL;
   output Vshamt;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   wire s_LOGISIM_NET_0;
   wire s_LOGISIM_NET_1;
   wire s_LOGISIM_NET_10;
   wire s_LOGISIM_NET_100;
   wire s_LOGISIM_NET_101;
   wire s_LOGISIM_NET_102;
   wire s_LOGISIM_NET_103;
   wire s_LOGISIM_NET_104;
   wire s_LOGISIM_NET_105;
   wire s_LOGISIM_NET_106;
   wire s_LOGISIM_NET_107;
   wire s_LOGISIM_NET_108;
   wire s_LOGISIM_NET_109;
   wire s_LOGISIM_NET_11;
   wire s_LOGISIM_NET_110;
   wire s_LOGISIM_NET_111;
   wire s_LOGISIM_NET_112;
   wire s_LOGISIM_NET_113;
   wire s_LOGISIM_NET_114;
   wire s_LOGISIM_NET_115;
   wire s_LOGISIM_NET_116;
   wire s_LOGISIM_NET_117;
   wire s_LOGISIM_NET_118;
   wire s_LOGISIM_NET_119;
   wire s_LOGISIM_NET_12;
   wire s_LOGISIM_NET_120;
   wire s_LOGISIM_NET_121;
   wire s_LOGISIM_NET_122;
   wire s_LOGISIM_NET_123;
   wire s_LOGISIM_NET_124;
   wire s_LOGISIM_NET_125;
   wire s_LOGISIM_NET_126;
   wire s_LOGISIM_NET_127;
   wire s_LOGISIM_NET_128;
   wire s_LOGISIM_NET_129;
   wire s_LOGISIM_NET_13;
   wire s_LOGISIM_NET_130;
   wire s_LOGISIM_NET_131;
   wire s_LOGISIM_NET_132;
   wire s_LOGISIM_NET_133;
   wire s_LOGISIM_NET_134;
   wire s_LOGISIM_NET_135;
   wire s_LOGISIM_NET_136;
   wire s_LOGISIM_NET_137;
   wire s_LOGISIM_NET_138;
   wire s_LOGISIM_NET_139;
   wire s_LOGISIM_NET_14;
   wire s_LOGISIM_NET_140;
   wire s_LOGISIM_NET_141;
   wire s_LOGISIM_NET_142;
   wire s_LOGISIM_NET_143;
   wire s_LOGISIM_NET_144;
   wire s_LOGISIM_NET_145;
   wire s_LOGISIM_NET_146;
   wire s_LOGISIM_NET_147;
   wire s_LOGISIM_NET_148;
   wire s_LOGISIM_NET_149;
   wire s_LOGISIM_NET_15;
   wire s_LOGISIM_NET_150;
   wire s_LOGISIM_NET_151;
   wire s_LOGISIM_NET_152;
   wire s_LOGISIM_NET_153;
   wire s_LOGISIM_NET_154;
   wire s_LOGISIM_NET_155;
   wire s_LOGISIM_NET_156;
   wire s_LOGISIM_NET_157;
   wire s_LOGISIM_NET_158;
   wire s_LOGISIM_NET_159;
   wire s_LOGISIM_NET_16;
   wire s_LOGISIM_NET_160;
   wire s_LOGISIM_NET_161;
   wire s_LOGISIM_NET_162;
   wire s_LOGISIM_NET_163;
   wire s_LOGISIM_NET_164;
   wire s_LOGISIM_NET_165;
   wire s_LOGISIM_NET_166;
   wire s_LOGISIM_NET_167;
   wire s_LOGISIM_NET_168;
   wire s_LOGISIM_NET_169;
   wire s_LOGISIM_NET_17;
   wire s_LOGISIM_NET_170;
   wire s_LOGISIM_NET_171;
   wire s_LOGISIM_NET_172;
   wire s_LOGISIM_NET_173;
   wire s_LOGISIM_NET_174;
   wire s_LOGISIM_NET_175;
   wire s_LOGISIM_NET_176;
   wire s_LOGISIM_NET_177;
   wire s_LOGISIM_NET_178;
   wire s_LOGISIM_NET_179;
   wire s_LOGISIM_NET_18;
   wire s_LOGISIM_NET_180;
   wire s_LOGISIM_NET_181;
   wire s_LOGISIM_NET_182;
   wire s_LOGISIM_NET_183;
   wire s_LOGISIM_NET_184;
   wire s_LOGISIM_NET_185;
   wire s_LOGISIM_NET_186;
   wire s_LOGISIM_NET_187;
   wire s_LOGISIM_NET_188;
   wire s_LOGISIM_NET_189;
   wire s_LOGISIM_NET_19;
   wire s_LOGISIM_NET_190;
   wire s_LOGISIM_NET_191;
   wire s_LOGISIM_NET_192;
   wire s_LOGISIM_NET_193;
   wire s_LOGISIM_NET_194;
   wire s_LOGISIM_NET_195;
   wire s_LOGISIM_NET_196;
   wire s_LOGISIM_NET_197;
   wire s_LOGISIM_NET_198;
   wire s_LOGISIM_NET_199;
   wire s_LOGISIM_NET_2;
   wire s_LOGISIM_NET_20;
   wire s_LOGISIM_NET_200;
   wire s_LOGISIM_NET_201;
   wire s_LOGISIM_NET_202;
   wire s_LOGISIM_NET_203;
   wire s_LOGISIM_NET_204;
   wire s_LOGISIM_NET_205;
   wire s_LOGISIM_NET_206;
   wire s_LOGISIM_NET_207;
   wire s_LOGISIM_NET_208;
   wire s_LOGISIM_NET_209;
   wire s_LOGISIM_NET_21;
   wire s_LOGISIM_NET_210;
   wire s_LOGISIM_NET_211;
   wire s_LOGISIM_NET_212;
   wire s_LOGISIM_NET_213;
   wire s_LOGISIM_NET_214;
   wire s_LOGISIM_NET_215;
   wire s_LOGISIM_NET_216;
   wire s_LOGISIM_NET_217;
   wire s_LOGISIM_NET_218;
   wire s_LOGISIM_NET_219;
   wire s_LOGISIM_NET_22;
   wire s_LOGISIM_NET_220;
   wire s_LOGISIM_NET_221;
   wire s_LOGISIM_NET_222;
   wire s_LOGISIM_NET_223;
   wire s_LOGISIM_NET_224;
   wire s_LOGISIM_NET_225;
   wire s_LOGISIM_NET_226;
   wire s_LOGISIM_NET_227;
   wire s_LOGISIM_NET_228;
   wire s_LOGISIM_NET_229;
   wire s_LOGISIM_NET_23;
   wire s_LOGISIM_NET_230;
   wire s_LOGISIM_NET_231;
   wire s_LOGISIM_NET_232;
   wire s_LOGISIM_NET_233;
   wire s_LOGISIM_NET_234;
   wire s_LOGISIM_NET_235;
   wire s_LOGISIM_NET_236;
   wire s_LOGISIM_NET_237;
   wire s_LOGISIM_NET_238;
   wire s_LOGISIM_NET_239;
   wire s_LOGISIM_NET_24;
   wire s_LOGISIM_NET_240;
   wire s_LOGISIM_NET_241;
   wire s_LOGISIM_NET_242;
   wire s_LOGISIM_NET_243;
   wire s_LOGISIM_NET_244;
   wire s_LOGISIM_NET_245;
   wire s_LOGISIM_NET_246;
   wire s_LOGISIM_NET_247;
   wire s_LOGISIM_NET_248;
   wire s_LOGISIM_NET_249;
   wire s_LOGISIM_NET_25;
   wire s_LOGISIM_NET_250;
   wire s_LOGISIM_NET_251;
   wire s_LOGISIM_NET_252;
   wire s_LOGISIM_NET_253;
   wire s_LOGISIM_NET_254;
   wire s_LOGISIM_NET_255;
   wire s_LOGISIM_NET_256;
   wire s_LOGISIM_NET_257;
   wire s_LOGISIM_NET_258;
   wire s_LOGISIM_NET_259;
   wire s_LOGISIM_NET_26;
   wire s_LOGISIM_NET_260;
   wire s_LOGISIM_NET_261;
   wire s_LOGISIM_NET_262;
   wire s_LOGISIM_NET_263;
   wire s_LOGISIM_NET_264;
   wire s_LOGISIM_NET_265;
   wire s_LOGISIM_NET_266;
   wire s_LOGISIM_NET_267;
   wire s_LOGISIM_NET_268;
   wire s_LOGISIM_NET_269;
   wire s_LOGISIM_NET_27;
   wire s_LOGISIM_NET_270;
   wire s_LOGISIM_NET_271;
   wire s_LOGISIM_NET_272;
   wire s_LOGISIM_NET_273;
   wire s_LOGISIM_NET_274;
   wire s_LOGISIM_NET_275;
   wire s_LOGISIM_NET_276;
   wire s_LOGISIM_NET_277;
   wire s_LOGISIM_NET_278;
   wire s_LOGISIM_NET_279;
   wire s_LOGISIM_NET_28;
   wire s_LOGISIM_NET_280;
   wire s_LOGISIM_NET_281;
   wire s_LOGISIM_NET_282;
   wire s_LOGISIM_NET_283;
   wire s_LOGISIM_NET_284;
   wire s_LOGISIM_NET_285;
   wire s_LOGISIM_NET_286;
   wire s_LOGISIM_NET_287;
   wire s_LOGISIM_NET_288;
   wire s_LOGISIM_NET_289;
   wire s_LOGISIM_NET_29;
   wire s_LOGISIM_NET_290;
   wire s_LOGISIM_NET_291;
   wire s_LOGISIM_NET_292;
   wire s_LOGISIM_NET_293;
   wire s_LOGISIM_NET_294;
   wire s_LOGISIM_NET_295;
   wire s_LOGISIM_NET_296;
   wire s_LOGISIM_NET_297;
   wire s_LOGISIM_NET_298;
   wire s_LOGISIM_NET_299;
   wire s_LOGISIM_NET_3;
   wire s_LOGISIM_NET_30;
   wire s_LOGISIM_NET_300;
   wire s_LOGISIM_NET_301;
   wire s_LOGISIM_NET_302;
   wire s_LOGISIM_NET_303;
   wire s_LOGISIM_NET_304;
   wire s_LOGISIM_NET_305;
   wire s_LOGISIM_NET_306;
   wire s_LOGISIM_NET_307;
   wire s_LOGISIM_NET_308;
   wire s_LOGISIM_NET_309;
   wire s_LOGISIM_NET_31;
   wire s_LOGISIM_NET_310;
   wire s_LOGISIM_NET_311;
   wire s_LOGISIM_NET_312;
   wire s_LOGISIM_NET_313;
   wire s_LOGISIM_NET_314;
   wire s_LOGISIM_NET_315;
   wire s_LOGISIM_NET_316;
   wire s_LOGISIM_NET_317;
   wire s_LOGISIM_NET_318;
   wire s_LOGISIM_NET_319;
   wire s_LOGISIM_NET_32;
   wire s_LOGISIM_NET_320;
   wire s_LOGISIM_NET_321;
   wire s_LOGISIM_NET_322;
   wire s_LOGISIM_NET_323;
   wire s_LOGISIM_NET_324;
   wire s_LOGISIM_NET_325;
   wire s_LOGISIM_NET_326;
   wire s_LOGISIM_NET_327;
   wire s_LOGISIM_NET_328;
   wire s_LOGISIM_NET_329;
   wire s_LOGISIM_NET_33;
   wire s_LOGISIM_NET_330;
   wire s_LOGISIM_NET_331;
   wire s_LOGISIM_NET_332;
   wire s_LOGISIM_NET_333;
   wire s_LOGISIM_NET_334;
   wire s_LOGISIM_NET_335;
   wire s_LOGISIM_NET_336;
   wire s_LOGISIM_NET_337;
   wire s_LOGISIM_NET_338;
   wire s_LOGISIM_NET_339;
   wire s_LOGISIM_NET_34;
   wire s_LOGISIM_NET_340;
   wire s_LOGISIM_NET_341;
   wire s_LOGISIM_NET_342;
   wire s_LOGISIM_NET_343;
   wire s_LOGISIM_NET_344;
   wire s_LOGISIM_NET_345;
   wire s_LOGISIM_NET_346;
   wire s_LOGISIM_NET_347;
   wire s_LOGISIM_NET_348;
   wire s_LOGISIM_NET_349;
   wire s_LOGISIM_NET_35;
   wire s_LOGISIM_NET_350;
   wire s_LOGISIM_NET_351;
   wire s_LOGISIM_NET_352;
   wire s_LOGISIM_NET_353;
   wire s_LOGISIM_NET_354;
   wire s_LOGISIM_NET_355;
   wire s_LOGISIM_NET_356;
   wire s_LOGISIM_NET_357;
   wire s_LOGISIM_NET_358;
   wire s_LOGISIM_NET_359;
   wire s_LOGISIM_NET_36;
   wire s_LOGISIM_NET_360;
   wire s_LOGISIM_NET_361;
   wire s_LOGISIM_NET_362;
   wire s_LOGISIM_NET_363;
   wire s_LOGISIM_NET_364;
   wire s_LOGISIM_NET_365;
   wire s_LOGISIM_NET_366;
   wire s_LOGISIM_NET_367;
   wire s_LOGISIM_NET_368;
   wire s_LOGISIM_NET_369;
   wire s_LOGISIM_NET_37;
   wire s_LOGISIM_NET_370;
   wire s_LOGISIM_NET_371;
   wire s_LOGISIM_NET_372;
   wire s_LOGISIM_NET_373;
   wire s_LOGISIM_NET_374;
   wire s_LOGISIM_NET_375;
   wire s_LOGISIM_NET_376;
   wire s_LOGISIM_NET_377;
   wire s_LOGISIM_NET_378;
   wire s_LOGISIM_NET_379;
   wire s_LOGISIM_NET_38;
   wire s_LOGISIM_NET_380;
   wire s_LOGISIM_NET_381;
   wire s_LOGISIM_NET_382;
   wire s_LOGISIM_NET_383;
   wire s_LOGISIM_NET_384;
   wire s_LOGISIM_NET_385;
   wire s_LOGISIM_NET_386;
   wire s_LOGISIM_NET_387;
   wire s_LOGISIM_NET_388;
   wire s_LOGISIM_NET_389;
   wire s_LOGISIM_NET_39;
   wire s_LOGISIM_NET_390;
   wire s_LOGISIM_NET_391;
   wire s_LOGISIM_NET_392;
   wire s_LOGISIM_NET_393;
   wire s_LOGISIM_NET_394;
   wire s_LOGISIM_NET_395;
   wire s_LOGISIM_NET_396;
   wire s_LOGISIM_NET_397;
   wire s_LOGISIM_NET_398;
   wire s_LOGISIM_NET_399;
   wire s_LOGISIM_NET_4;
   wire s_LOGISIM_NET_40;
   wire s_LOGISIM_NET_400;
   wire s_LOGISIM_NET_401;
   wire s_LOGISIM_NET_402;
   wire s_LOGISIM_NET_403;
   wire s_LOGISIM_NET_404;
   wire s_LOGISIM_NET_405;
   wire s_LOGISIM_NET_406;
   wire s_LOGISIM_NET_407;
   wire s_LOGISIM_NET_408;
   wire s_LOGISIM_NET_409;
   wire s_LOGISIM_NET_41;
   wire s_LOGISIM_NET_410;
   wire s_LOGISIM_NET_411;
   wire s_LOGISIM_NET_412;
   wire s_LOGISIM_NET_413;
   wire s_LOGISIM_NET_414;
   wire s_LOGISIM_NET_415;
   wire s_LOGISIM_NET_416;
   wire s_LOGISIM_NET_417;
   wire s_LOGISIM_NET_418;
   wire s_LOGISIM_NET_419;
   wire s_LOGISIM_NET_42;
   wire s_LOGISIM_NET_420;
   wire s_LOGISIM_NET_421;
   wire s_LOGISIM_NET_422;
   wire s_LOGISIM_NET_423;
   wire s_LOGISIM_NET_424;
   wire s_LOGISIM_NET_425;
   wire s_LOGISIM_NET_426;
   wire s_LOGISIM_NET_427;
   wire s_LOGISIM_NET_428;
   wire s_LOGISIM_NET_429;
   wire s_LOGISIM_NET_43;
   wire s_LOGISIM_NET_430;
   wire s_LOGISIM_NET_431;
   wire s_LOGISIM_NET_432;
   wire s_LOGISIM_NET_433;
   wire s_LOGISIM_NET_434;
   wire s_LOGISIM_NET_435;
   wire s_LOGISIM_NET_436;
   wire s_LOGISIM_NET_437;
   wire s_LOGISIM_NET_438;
   wire s_LOGISIM_NET_439;
   wire s_LOGISIM_NET_44;
   wire s_LOGISIM_NET_440;
   wire s_LOGISIM_NET_441;
   wire s_LOGISIM_NET_442;
   wire s_LOGISIM_NET_443;
   wire s_LOGISIM_NET_444;
   wire s_LOGISIM_NET_445;
   wire s_LOGISIM_NET_446;
   wire s_LOGISIM_NET_447;
   wire s_LOGISIM_NET_448;
   wire s_LOGISIM_NET_449;
   wire s_LOGISIM_NET_45;
   wire s_LOGISIM_NET_450;
   wire s_LOGISIM_NET_451;
   wire s_LOGISIM_NET_452;
   wire s_LOGISIM_NET_453;
   wire s_LOGISIM_NET_454;
   wire s_LOGISIM_NET_455;
   wire s_LOGISIM_NET_456;
   wire s_LOGISIM_NET_457;
   wire s_LOGISIM_NET_458;
   wire s_LOGISIM_NET_459;
   wire s_LOGISIM_NET_46;
   wire s_LOGISIM_NET_460;
   wire s_LOGISIM_NET_461;
   wire s_LOGISIM_NET_462;
   wire s_LOGISIM_NET_463;
   wire s_LOGISIM_NET_464;
   wire s_LOGISIM_NET_465;
   wire s_LOGISIM_NET_466;
   wire s_LOGISIM_NET_467;
   wire s_LOGISIM_NET_468;
   wire s_LOGISIM_NET_469;
   wire s_LOGISIM_NET_47;
   wire s_LOGISIM_NET_470;
   wire s_LOGISIM_NET_471;
   wire s_LOGISIM_NET_472;
   wire s_LOGISIM_NET_473;
   wire s_LOGISIM_NET_474;
   wire s_LOGISIM_NET_475;
   wire s_LOGISIM_NET_476;
   wire s_LOGISIM_NET_477;
   wire s_LOGISIM_NET_478;
   wire s_LOGISIM_NET_479;
   wire s_LOGISIM_NET_48;
   wire s_LOGISIM_NET_480;
   wire s_LOGISIM_NET_49;
   wire s_LOGISIM_NET_5;
   wire s_LOGISIM_NET_50;
   wire s_LOGISIM_NET_51;
   wire s_LOGISIM_NET_52;
   wire s_LOGISIM_NET_53;
   wire s_LOGISIM_NET_54;
   wire s_LOGISIM_NET_55;
   wire s_LOGISIM_NET_56;
   wire s_LOGISIM_NET_57;
   wire s_LOGISIM_NET_58;
   wire s_LOGISIM_NET_59;
   wire s_LOGISIM_NET_6;
   wire s_LOGISIM_NET_60;
   wire s_LOGISIM_NET_61;
   wire s_LOGISIM_NET_62;
   wire s_LOGISIM_NET_63;
   wire s_LOGISIM_NET_64;
   wire s_LOGISIM_NET_65;
   wire s_LOGISIM_NET_66;
   wire s_LOGISIM_NET_67;
   wire s_LOGISIM_NET_68;
   wire s_LOGISIM_NET_69;
   wire s_LOGISIM_NET_7;
   wire s_LOGISIM_NET_70;
   wire s_LOGISIM_NET_71;
   wire s_LOGISIM_NET_72;
   wire s_LOGISIM_NET_73;
   wire s_LOGISIM_NET_74;
   wire s_LOGISIM_NET_75;
   wire s_LOGISIM_NET_76;
   wire s_LOGISIM_NET_77;
   wire s_LOGISIM_NET_78;
   wire s_LOGISIM_NET_79;
   wire s_LOGISIM_NET_8;
   wire s_LOGISIM_NET_80;
   wire s_LOGISIM_NET_81;
   wire s_LOGISIM_NET_82;
   wire s_LOGISIM_NET_83;
   wire s_LOGISIM_NET_84;
   wire s_LOGISIM_NET_85;
   wire s_LOGISIM_NET_86;
   wire s_LOGISIM_NET_87;
   wire s_LOGISIM_NET_88;
   wire s_LOGISIM_NET_89;
   wire s_LOGISIM_NET_9;
   wire s_LOGISIM_NET_90;
   wire s_LOGISIM_NET_91;
   wire s_LOGISIM_NET_92;
   wire s_LOGISIM_NET_93;
   wire s_LOGISIM_NET_94;
   wire s_LOGISIM_NET_95;
   wire s_LOGISIM_NET_96;
   wire s_LOGISIM_NET_97;
   wire s_LOGISIM_NET_98;
   wire s_LOGISIM_NET_99;


   /***************************************************************************
    ** Here all input connections are defined                                **
    ***************************************************************************/
   assign s_LOGISIM_NET_42                   = F4;
   assign s_LOGISIM_NET_30                   = F2;
   assign s_LOGISIM_NET_5                    = OP4;
   assign s_LOGISIM_NET_27                   = OP3;
   assign s_LOGISIM_NET_10                   = F1;
   assign s_LOGISIM_NET_37                   = OP0;
   assign s_LOGISIM_NET_14                   = F0;
   assign s_LOGISIM_NET_6                    = OP5;
   assign s_LOGISIM_NET_88                   = F3;
   assign s_LOGISIM_NET_11                   = OP2;
   assign s_LOGISIM_NET_12                   = OP1;
   assign s_LOGISIM_NET_7                    = F5;

   /***************************************************************************
    ** Here all output connections are defined                               **
    ***************************************************************************/
   assign MemToReg                           = s_LOGISIM_NET_361;
   assign SignedExt                          = s_LOGISIM_NET_284;
   assign JUMP                               = s_LOGISIM_NET_445;
   assign RegDst                             = s_LOGISIM_NET_163;
   assign BNE                                = s_LOGISIM_NET_475;
   assign Vshamt                             = s_LOGISIM_NET_463;
   assign SysCALL                            = s_LOGISIM_NET_426;
   assign MemWrite                           = s_LOGISIM_NET_126;
   assign JAL                                = s_LOGISIM_NET_476;
   assign BLEZ                               = s_LOGISIM_NET_381;
   assign BEQ                                = s_LOGISIM_NET_444;
   assign JR                                 = s_LOGISIM_NET_462;
   assign HalfW                              = s_LOGISIM_NET_431;
   assign RegWrite                           = s_LOGISIM_NET_413;
   assign ALU_SRC                            = s_LOGISIM_NET_241;

   /***************************************************************************
    ** Here all normal components are defined                                **
    ***************************************************************************/
   NOT_GATE      GATE_1 (.Input_1(s_LOGISIM_NET_27),
                         .Result(s_LOGISIM_NET_457));

   NOT_GATE      GATE_2 (.Input_1(s_LOGISIM_NET_11),
                         .Result(s_LOGISIM_NET_465));

   NOT_GATE      GATE_3 (.Input_1(s_LOGISIM_NET_27),
                         .Result(s_LOGISIM_NET_379));

   NOT_GATE      GATE_4 (.Input_1(s_LOGISIM_NET_37),
                         .Result(s_LOGISIM_NET_478));

   NOT_GATE      GATE_5 (.Input_1(s_LOGISIM_NET_37),
                         .Result(s_LOGISIM_NET_461));

   NOT_GATE      GATE_6 (.Input_1(s_LOGISIM_NET_6),
                         .Result(s_LOGISIM_NET_164));

   NOT_GATE      GATE_7 (.Input_1(s_LOGISIM_NET_37),
                         .Result(s_LOGISIM_NET_8));

   NOT_GATE      GATE_8 (.Input_1(s_LOGISIM_NET_5),
                         .Result(s_LOGISIM_NET_136));

   NOT_GATE      GATE_9 (.Input_1(s_LOGISIM_NET_12),
                         .Result(s_LOGISIM_NET_443));

   NOT_GATE      GATE_10 (.Input_1(s_LOGISIM_NET_11),
                          .Result(s_LOGISIM_NET_177));

   NOT_GATE      GATE_11 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_234));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_12 (.Input_1(s_LOGISIM_NET_6),
               .Input_2(s_LOGISIM_NET_220),
               .Input_3(s_LOGISIM_NET_27),
               .Input_4(s_LOGISIM_NET_454),
               .Input_5(s_LOGISIM_NET_430),
               .Input_6(s_LOGISIM_NET_37),
               .Result(s_LOGISIM_NET_342));

   NOT_GATE      GATE_13 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_264));

   NOT_GATE      GATE_14 (.Input_1(s_LOGISIM_NET_88),
                          .Result(s_LOGISIM_NET_295));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_15 (.Input_1(s_LOGISIM_NET_37),
               .Input_2(s_LOGISIM_NET_192),
               .Input_3(s_LOGISIM_NET_429),
               .Input_4(s_LOGISIM_NET_27),
               .Input_5(s_LOGISIM_NET_436),
               .Input_6(s_LOGISIM_NET_6),
               .Result(s_LOGISIM_NET_431));

   NOT_GATE      GATE_16 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_337));

   NOT_GATE      GATE_17 (.Input_1(s_LOGISIM_NET_27),
                          .Result(s_LOGISIM_NET_195));

   NOT_GATE      GATE_18 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_168));

   NOT_GATE      GATE_19 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_406));

   NOT_GATE      GATE_20 (.Input_1(s_LOGISIM_NET_10),
                          .Result(s_LOGISIM_NET_213));

   NOT_GATE      GATE_21 (.Input_1(s_LOGISIM_NET_11),
                          .Result(s_LOGISIM_NET_259));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_22 (.Input_1(s_LOGISIM_NET_62),
               .Input_10(s_LOGISIM_NET_152),
               .Input_11(s_LOGISIM_NET_319),
               .Input_12(s_LOGISIM_NET_14),
               .Input_2(s_LOGISIM_NET_458),
               .Input_3(s_LOGISIM_NET_3),
               .Input_4(s_LOGISIM_NET_177),
               .Input_5(s_LOGISIM_NET_309),
               .Input_6(s_LOGISIM_NET_18),
               .Input_7(s_LOGISIM_NET_7),
               .Input_8(s_LOGISIM_NET_277),
               .Input_9(s_LOGISIM_NET_184),
               .Result(s_LOGISIM_NET_420));

   NOT_GATE      GATE_23 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_334));

   NOT_GATE      GATE_24 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_63));

   NOT_GATE      GATE_25 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_346));

   NOT_GATE      GATE_26 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_23));

   NOT_GATE      GATE_27 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_375));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_28 (.Input_1(s_LOGISIM_NET_385),
               .Input_10(s_LOGISIM_NET_30),
               .Input_11(s_LOGISIM_NET_173),
               .Input_12(s_LOGISIM_NET_433),
               .Input_2(s_LOGISIM_NET_415),
               .Input_3(s_LOGISIM_NET_307),
               .Input_4(s_LOGISIM_NET_68),
               .Input_5(s_LOGISIM_NET_159),
               .Input_6(s_LOGISIM_NET_466),
               .Input_7(s_LOGISIM_NET_162),
               .Input_8(s_LOGISIM_NET_113),
               .Input_9(s_LOGISIM_NET_88),
               .Result(s_LOGISIM_NET_426));

   NOT_GATE      GATE_29 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_414));

   NOT_GATE      GATE_30 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_64));

   NOT_GATE      GATE_31 (.Input_1(s_LOGISIM_NET_27),
                          .Result(s_LOGISIM_NET_307));

   NOT_GATE      GATE_32 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_108));

   NOT_GATE      GATE_33 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_36));

   NOT_GATE      GATE_34 (.Input_1(s_LOGISIM_NET_88),
                          .Result(s_LOGISIM_NET_101));

   NOT_GATE      GATE_35 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_385));

   NOT_GATE      GATE_36 (.Input_1(s_LOGISIM_NET_27),
                          .Result(s_LOGISIM_NET_111));

   NOT_GATE      GATE_37 (.Input_1(s_LOGISIM_NET_42),
                          .Result(s_LOGISIM_NET_392));

   NOT_GATE      GATE_38 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_123));

   NOT_GATE      GATE_39 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_94));

   NOT_GATE      GATE_40 (.Input_1(s_LOGISIM_NET_37),
                          .Result(s_LOGISIM_NET_351));

   NOT_GATE      GATE_41 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_286));

   NOT_GATE      GATE_42 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_453));

   NOT_GATE      GATE_43 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_451));

   NOT_GATE      GATE_44 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_355));

   NOT_GATE      GATE_45 (.Input_1(s_LOGISIM_NET_11),
                          .Result(s_LOGISIM_NET_370));

   NOT_GATE      GATE_46 (.Input_1(s_LOGISIM_NET_88),
                          .Result(s_LOGISIM_NET_133));

   NOT_GATE      GATE_47 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_291));

   NOT_GATE      GATE_48 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_382));

   NOT_GATE      GATE_49 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_102));

   NOT_GATE      GATE_50 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_327));

   NOT_GATE      GATE_51 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_464));

   NOT_GATE      GATE_52 (.Input_1(s_LOGISIM_NET_42),
                          .Result(s_LOGISIM_NET_40));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_53 (.Input_1(s_LOGISIM_NET_36),
               .Input_2(s_LOGISIM_NET_193),
               .Input_3(s_LOGISIM_NET_427),
               .Input_4(s_LOGISIM_NET_11),
               .Input_5(s_LOGISIM_NET_437),
               .Input_6(s_LOGISIM_NET_37),
               .Result(s_LOGISIM_NET_280));

   NOT_GATE      GATE_54 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_110));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_55 (.Input_1(s_LOGISIM_NET_180),
               .Input_2(s_LOGISIM_NET_327),
               .Input_3(s_LOGISIM_NET_343),
               .Input_4(s_LOGISIM_NET_11),
               .Input_5(s_LOGISIM_NET_366),
               .Input_6(s_LOGISIM_NET_106),
               .Result(s_LOGISIM_NET_186));

   NOT_GATE      GATE_56 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_200));

   NOT_GATE      GATE_57 (.Input_1(s_LOGISIM_NET_27),
                          .Result(s_LOGISIM_NET_143));

   NOT_GATE      GATE_58 (.Input_1(s_LOGISIM_NET_27),
                          .Result(s_LOGISIM_NET_253));

   NOT_GATE      GATE_59 (.Input_1(s_LOGISIM_NET_88),
                          .Result(s_LOGISIM_NET_403));

   NOT_GATE      GATE_60 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_417));

   NOT_GATE      GATE_61 (.Input_1(s_LOGISIM_NET_11),
                          .Result(s_LOGISIM_NET_97));

   NOT_GATE      GATE_62 (.Input_1(s_LOGISIM_NET_37),
                          .Result(s_LOGISIM_NET_265));

   NOT_GATE      GATE_63 (.Input_1(s_LOGISIM_NET_37),
                          .Result(s_LOGISIM_NET_339));

   NOT_GATE      GATE_64 (.Input_1(s_LOGISIM_NET_30),
                          .Result(s_LOGISIM_NET_51));

   NOT_GATE      GATE_65 (.Input_1(s_LOGISIM_NET_27),
                          .Result(s_LOGISIM_NET_474));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_66 (.Input_1(s_LOGISIM_NET_77),
               .Input_10(s_LOGISIM_NET_33),
               .Input_11(s_LOGISIM_NET_311),
               .Input_12(s_LOGISIM_NET_231),
               .Input_2(s_LOGISIM_NET_167),
               .Input_3(s_LOGISIM_NET_142),
               .Input_4(s_LOGISIM_NET_399),
               .Input_5(s_LOGISIM_NET_321),
               .Input_6(s_LOGISIM_NET_340),
               .Input_7(s_LOGISIM_NET_108),
               .Input_8(s_LOGISIM_NET_217),
               .Input_9(s_LOGISIM_NET_99),
               .Result(s_LOGISIM_NET_214));

   NOT_GATE      GATE_67 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_219));

   NOT_GATE      GATE_68 (.Input_1(s_LOGISIM_NET_11),
                          .Result(s_LOGISIM_NET_146));

   NOT_GATE      GATE_69 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_77));

   NOT_GATE      GATE_70 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_424));

   NOT_GATE      GATE_71 (.Input_1(s_LOGISIM_NET_27),
                          .Result(s_LOGISIM_NET_3));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_72 (.Input_1(s_LOGISIM_NET_188),
               .Input_2(s_LOGISIM_NET_382),
               .Input_3(s_LOGISIM_NET_473),
               .Input_4(s_LOGISIM_NET_11),
               .Input_5(s_LOGISIM_NET_0),
               .Input_6(s_LOGISIM_NET_37),
               .Result(s_LOGISIM_NET_475));

   NOT_GATE      GATE_73 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_331));

   NOT_GATE      GATE_74 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_155));

   NOT_GATE      GATE_75 (.Input_1(s_LOGISIM_NET_27),
                          .Result(s_LOGISIM_NET_115));

   OR_GATE_20_INPUTS #(.BubblesMask(0))
      GATE_76 (.Input_1(s_LOGISIM_NET_214),
               .Input_10(s_LOGISIM_NET_270),
               .Input_11(s_LOGISIM_NET_360),
               .Input_12(s_LOGISIM_NET_182),
               .Input_13(s_LOGISIM_NET_275),
               .Input_14(s_LOGISIM_NET_238),
               .Input_15(s_LOGISIM_NET_141),
               .Input_16(s_LOGISIM_NET_297),
               .Input_17(s_LOGISIM_NET_407),
               .Input_18(s_LOGISIM_NET_329),
               .Input_19(s_LOGISIM_NET_367),
               .Input_2(s_LOGISIM_NET_350),
               .Input_20(s_LOGISIM_NET_243),
               .Input_3(s_LOGISIM_NET_165),
               .Input_4(s_LOGISIM_NET_353),
               .Input_5(s_LOGISIM_NET_420),
               .Input_6(s_LOGISIM_NET_316),
               .Input_7(s_LOGISIM_NET_95),
               .Input_8(s_LOGISIM_NET_268),
               .Input_9(s_LOGISIM_NET_398),
               .Result(s_LOGISIM_NET_413));

   NOT_GATE      GATE_77 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_404));

   NOT_GATE      GATE_78 (.Input_1(s_LOGISIM_NET_37),
                          .Result(s_LOGISIM_NET_59));

   NOT_GATE      GATE_79 (.Input_1(s_LOGISIM_NET_11),
                          .Result(s_LOGISIM_NET_85));

   NOT_GATE      GATE_80 (.Input_1(s_LOGISIM_NET_30),
                          .Result(s_LOGISIM_NET_239));

   NOT_GATE      GATE_81 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_39));

   NOT_GATE      GATE_82 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_289));

   NOT_GATE      GATE_83 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_368));

   NOT_GATE      GATE_84 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_371));

   NOT_GATE      GATE_85 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_363));

   NOT_GATE      GATE_86 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_421));

   NOT_GATE      GATE_87 (.Input_1(s_LOGISIM_NET_42),
                          .Result(s_LOGISIM_NET_139));

   NOT_GATE      GATE_88 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_89));

   NOT_GATE      GATE_89 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_292));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_90 (.Input_1(s_LOGISIM_NET_64),
               .Input_10(s_LOGISIM_NET_56),
               .Input_11(s_LOGISIM_NET_10),
               .Input_12(s_LOGISIM_NET_455),
               .Input_2(s_LOGISIM_NET_434),
               .Input_3(s_LOGISIM_NET_347),
               .Input_4(s_LOGISIM_NET_83),
               .Input_5(s_LOGISIM_NET_234),
               .Input_6(s_LOGISIM_NET_472),
               .Input_7(s_LOGISIM_NET_7),
               .Input_8(s_LOGISIM_NET_201),
               .Input_9(s_LOGISIM_NET_100),
               .Result(s_LOGISIM_NET_262));

   NOT_GATE      GATE_91 (.Input_1(s_LOGISIM_NET_11),
                          .Result(s_LOGISIM_NET_75));

   NOT_GATE      GATE_92 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_276));

   NOT_GATE      GATE_93 (.Input_1(s_LOGISIM_NET_5),
                          .Result(s_LOGISIM_NET_422));

   NOT_GATE      GATE_94 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_87));

   NOT_GATE      GATE_95 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_153));

   NOT_GATE      GATE_96 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_107));

   NOT_GATE      GATE_97 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_287));

   NOT_GATE      GATE_98 (.Input_1(s_LOGISIM_NET_6),
                          .Result(s_LOGISIM_NET_76));

   NOT_GATE      GATE_99 (.Input_1(s_LOGISIM_NET_11),
                          .Result(s_LOGISIM_NET_386));

   NOT_GATE      GATE_100 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_347));

   NOT_GATE      GATE_101 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_246));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_102 (.Input_1(s_LOGISIM_NET_63),
                .Input_10(s_LOGISIM_NET_30),
                .Input_11(s_LOGISIM_NET_318),
                .Input_12(s_LOGISIM_NET_468),
                .Input_2(s_LOGISIM_NET_459),
                .Input_3(s_LOGISIM_NET_4),
                .Input_4(s_LOGISIM_NET_178),
                .Input_5(s_LOGISIM_NET_310),
                .Input_6(s_LOGISIM_NET_19),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_279),
                .Input_9(s_LOGISIM_NET_185),
                .Result(s_LOGISIM_NET_95));

   NOT_GATE      GATE_103 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_383));

   NOT_GATE      GATE_104 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_120));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_105 (.Input_1(s_LOGISIM_NET_76),
                .Input_10(s_LOGISIM_NET_216),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_169),
                .Input_3(s_LOGISIM_NET_143),
                .Input_4(s_LOGISIM_NET_401),
                .Input_5(s_LOGISIM_NET_322),
                .Input_6(s_LOGISIM_NET_339),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_212),
                .Input_9(s_LOGISIM_NET_88),
                .Result(s_LOGISIM_NET_360));

   NOT_GATE      GATE_106 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_251));

   NOT_GATE      GATE_107 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_305));

   NOT_GATE      GATE_108 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_34));

   NOT_GATE      GATE_109 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_175));

   NOT_GATE      GATE_110 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_412));

   NOT_GATE      GATE_111 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_24));

   NOT_GATE      GATE_112 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_169));

   NOT_GATE      GATE_113 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_306));

   NOT_GATE      GATE_114 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_134));

   NOT_GATE      GATE_115 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_22));

   NOT_GATE      GATE_116 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_196));

   NOT_GATE      GATE_117 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_233));

   NOT_GATE      GATE_118 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_181));

   NOT_GATE      GATE_119 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_13));

   NOT_GATE      GATE_120 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_479));

   NOT_GATE      GATE_121 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_56));

   NOT_GATE      GATE_122 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_173));

   NOT_GATE      GATE_123 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_26));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_124 (.Input_1(s_LOGISIM_NET_196),
                .Input_10(s_LOGISIM_NET_317),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_320),
                .Input_2(s_LOGISIM_NET_272),
                .Input_3(s_LOGISIM_NET_17),
                .Input_4(s_LOGISIM_NET_74),
                .Input_5(s_LOGISIM_NET_375),
                .Input_6(s_LOGISIM_NET_389),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_313),
                .Input_9(s_LOGISIM_NET_210),
                .Result(s_LOGISIM_NET_316));

   NOT_GATE      GATE_125 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_116));

   NOT_GATE      GATE_126 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_192));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_127 (.Input_1(s_LOGISIM_NET_140),
                .Input_10(s_LOGISIM_NET_269),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_235),
                .Input_2(s_LOGISIM_NET_219),
                .Input_3(s_LOGISIM_NET_195),
                .Input_4(s_LOGISIM_NET_418),
                .Input_5(s_LOGISIM_NET_346),
                .Input_6(s_LOGISIM_NET_369),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_266),
                .Input_9(s_LOGISIM_NET_88),
                .Result(s_LOGISIM_NET_278));

   NOT_GATE      GATE_128 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_281));

   NOT_GATE      GATE_129 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_58));

   NOT_GATE      GATE_130 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_80));

   NOT_GATE      GATE_131 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_380));

   NOT_GATE      GATE_132 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_458));

   NOT_GATE      GATE_133 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_345));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_134 (.Input_1(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_187),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_447),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_218));

   NOT_GATE      GATE_135 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_387));

   NOT_GATE      GATE_136 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_69));

   NOT_GATE      GATE_137 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_271));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_138 (.Input_1(s_LOGISIM_NET_373),
                .Input_10(s_LOGISIM_NET_130),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_404),
                .Input_3(s_LOGISIM_NET_282),
                .Input_4(s_LOGISIM_NET_31),
                .Input_5(s_LOGISIM_NET_120),
                .Input_6(s_LOGISIM_NET_460),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_82),
                .Input_9(s_LOGISIM_NET_88),
                .Result(s_LOGISIM_NET_440));

   NOT_GATE      GATE_139 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_193));

   NOT_GATE      GATE_140 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_232));

   NOT_GATE      GATE_141 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_310));

   NOT_GATE      GATE_142 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_184));

   NOT_GATE      GATE_143 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_330));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_144 (.Input_1(s_LOGISIM_NET_20),
                .Input_10(s_LOGISIM_NET_30),
                .Input_11(s_LOGISIM_NET_304),
                .Input_12(s_LOGISIM_NET_93),
                .Input_2(s_LOGISIM_NET_452),
                .Input_3(s_LOGISIM_NET_380),
                .Input_4(s_LOGISIM_NET_149),
                .Input_5(s_LOGISIM_NET_289),
                .Input_6(s_LOGISIM_NET_480),
                .Input_7(s_LOGISIM_NET_292),
                .Input_8(s_LOGISIM_NET_258),
                .Input_9(s_LOGISIM_NET_296),
                .Result(s_LOGISIM_NET_463));

   NOT_GATE      GATE_145 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_45));

   NOT_GATE      GATE_146 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_466));

   NOT_GATE      GATE_147 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_43));

   NOT_GATE      GATE_148 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_159));

   NOT_GATE      GATE_149 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_237));

   NOT_GATE      GATE_150 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_180));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_151 (.Input_1(s_LOGISIM_NET_23),
                .Input_10(s_LOGISIM_NET_30),
                .Input_11(s_LOGISIM_NET_305),
                .Input_12(s_LOGISIM_NET_91),
                .Input_2(s_LOGISIM_NET_450),
                .Input_3(s_LOGISIM_NET_378),
                .Input_4(s_LOGISIM_NET_146),
                .Input_5(s_LOGISIM_NET_287),
                .Input_6(s_LOGISIM_NET_478),
                .Input_7(s_LOGISIM_NET_290),
                .Input_8(s_LOGISIM_NET_256),
                .Input_9(s_LOGISIM_NET_295),
                .Result(s_LOGISIM_NET_207));

   NOT_GATE      GATE_152 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_50));

   NOT_GATE      GATE_153 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_319));

   NOT_GATE      GATE_154 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_396));

   NOT_GATE      GATE_155 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_73));

   NOT_GATE      GATE_156 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_411));

   NOT_GATE      GATE_157 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_376));

   NOT_GATE      GATE_158 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_369));

   NOT_GATE      GATE_159 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_244));

   NOT_GATE      GATE_160 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_0));

   NOT_GATE      GATE_161 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_245));

   NOT_GATE      GATE_162 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_190));

   NOT_GATE      GATE_163 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_395));

   NOT_GATE      GATE_164 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_349));

   NOT_GATE      GATE_165 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_74));

   NOT_GATE      GATE_166 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_142));

   NOT_GATE      GATE_167 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_303));

   NOT_GATE      GATE_168 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_279));

   NOT_GATE      GATE_169 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_447));

   NOT_GATE      GATE_170 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_301));

   NOT_GATE      GATE_171 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_212));

   NOT_GATE      GATE_172 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_79));

   NOT_GATE      GATE_173 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_103));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_174 (.Input_1(s_LOGISIM_NET_103),
                .Input_2(s_LOGISIM_NET_247),
                .Input_3(s_LOGISIM_NET_442),
                .Input_4(s_LOGISIM_NET_252),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_118),
                .Result(s_LOGISIM_NET_445));

   NOT_GATE      GATE_175 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_344));

   NOT_GATE      GATE_176 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_389));

   NOT_GATE      GATE_177 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_152));

   NOT_GATE      GATE_178 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_325));

   NOT_GATE      GATE_179 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_154));

   NOT_GATE      GATE_180 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_419));

   NOT_GATE      GATE_181 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_269));

   NOT_GATE      GATE_182 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_338));

   NOT_GATE      GATE_183 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_66));

   NOT_GATE      GATE_184 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_441));

   NOT_GATE      GATE_185 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_137));

   NOT_GATE      GATE_186 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_226));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_187 (.Input_1(s_LOGISIM_NET_276),
                .Input_10(s_LOGISIM_NET_239),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_331),
                .Input_3(s_LOGISIM_NET_115),
                .Input_4(s_LOGISIM_NET_166),
                .Input_5(s_LOGISIM_NET_409),
                .Input_6(s_LOGISIM_NET_419),
                .Input_7(s_LOGISIM_NET_299),
                .Input_8(s_LOGISIM_NET_359),
                .Input_9(s_LOGISIM_NET_293),
                .Result(s_LOGISIM_NET_391));

   NOT_GATE      GATE_188 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_252));

   NOT_GATE      GATE_189 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_203));

   NOT_GATE      GATE_190 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_277));

   NOT_GATE      GATE_191 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_373));

   NOT_GATE      GATE_192 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_358));

   NOT_GATE      GATE_193 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_254));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_194 (.Input_1(s_LOGISIM_NET_60),
                .Input_2(s_LOGISIM_NET_362),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_477),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_135));

   NOT_GATE      GATE_195 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_437));

   NOT_GATE      GATE_196 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_84));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_197 (.Input_1(s_LOGISIM_NET_39),
                .Input_2(s_LOGISIM_NET_158),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_11),
                .Input_5(s_LOGISIM_NET_222),
                .Input_6(s_LOGISIM_NET_412),
                .Result(s_LOGISIM_NET_238));

   NOT_GATE      GATE_198 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_242));

   NOT_GATE      GATE_199 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_52));

   NOT_GATE      GATE_200 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_477));

   NOT_GATE      GATE_201 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_220));

   NOT_GATE      GATE_202 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_272));

   NOT_GATE      GATE_203 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_71));

   NOT_GATE      GATE_204 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_202));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_205 (.Input_1(s_LOGISIM_NET_102),
                .Input_2(s_LOGISIM_NET_246),
                .Input_3(s_LOGISIM_NET_441),
                .Input_4(s_LOGISIM_NET_11),
                .Input_5(s_LOGISIM_NET_453),
                .Input_6(s_LOGISIM_NET_116),
                .Result(s_LOGISIM_NET_444));

   NOT_GATE      GATE_206 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_348));

   NOT_GATE      GATE_207 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_149));

   NOT_GATE      GATE_208 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_127));

   NOT_GATE      GATE_209 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_191));

   NOT_GATE      GATE_210 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_15));

   NOT_GATE      GATE_211 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_187));

   NOT_GATE      GATE_212 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_317));

   NOT_GATE      GATE_213 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_46));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_214 (.Input_1(s_LOGISIM_NET_156),
                .Input_10(s_LOGISIM_NET_226),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_87),
                .Input_2(s_LOGISIM_NET_57),
                .Input_3(s_LOGISIM_NET_112),
                .Input_4(s_LOGISIM_NET_259),
                .Input_5(s_LOGISIM_NET_81),
                .Input_6(s_LOGISIM_NET_125),
                .Input_7(s_LOGISIM_NET_355),
                .Input_8(s_LOGISIM_NET_139),
                .Input_9(s_LOGISIM_NET_357),
                .Result(s_LOGISIM_NET_448));

   NOT_GATE      GATE_215 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_176));

   NOT_GATE      GATE_216 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_235));

   NOT_GATE      GATE_217 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_455));

   NOT_GATE      GATE_218 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_410));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_219 (.Input_1(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_9),
                .Input_3(s_LOGISIM_NET_354),
                .Input_4(s_LOGISIM_NET_271),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_361));

   NOT_GATE      GATE_220 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_399));

   NOT_GATE      GATE_221 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_427));

   NOT_GATE      GATE_222 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_230));

   NOT_GATE      GATE_223 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_32));

   NOT_GATE      GATE_224 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_201));

   NOT_GATE      GATE_225 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_249));

   NOT_GATE      GATE_226 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_432));

   NOT_GATE      GATE_227 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_274));

   NOT_GATE      GATE_228 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_282));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_229 (.Input_1(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_244),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_364),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_25));

   NOT_GATE      GATE_230 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_17));

   NOT_GATE      GATE_231 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_86));

   NOT_GATE      GATE_232 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_288));

   OR_GATE #(.BubblesMask(0))
      GATE_233 (.Input_1(s_LOGISIM_NET_25),
                .Input_2(s_LOGISIM_NET_49),
                .Result(s_LOGISIM_NET_126));

   NOT_GATE      GATE_234 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_312));

   NOT_GATE      GATE_235 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_313));

   NOT_GATE      GATE_236 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_185));

   NOT_GATE      GATE_237 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_55));

   NOT_GATE      GATE_238 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_128));

   NOT_GATE      GATE_239 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_183));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_240 (.Input_1(s_LOGISIM_NET_109),
                .Input_10(s_LOGISIM_NET_250),
                .Input_11(s_LOGISIM_NET_213),
                .Input_12(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_190),
                .Input_3(s_LOGISIM_NET_171),
                .Input_4(s_LOGISIM_NET_410),
                .Input_5(s_LOGISIM_NET_334),
                .Input_6(s_LOGISIM_NET_351),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_236),
                .Input_9(s_LOGISIM_NET_128),
                .Result(s_LOGISIM_NET_122));

   NOT_GATE      GATE_241 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_359));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_242 (.Input_1(s_LOGISIM_NET_153),
                .Input_2(s_LOGISIM_NET_368),
                .Input_3(s_LOGISIM_NET_470),
                .Input_4(s_LOGISIM_NET_370),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_182));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_243 (.Input_1(s_LOGISIM_NET_261),
                .Input_2(s_LOGISIM_NET_46),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_11),
                .Input_5(s_LOGISIM_NET_371),
                .Input_6(s_LOGISIM_NET_121),
                .Result(s_LOGISIM_NET_151));

   NOT_GATE      GATE_244 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_356));

   NOT_GATE      GATE_245 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_418));

   NOT_GATE      GATE_246 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_460));

   NOT_GATE      GATE_247 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_16));

   NOT_GATE      GATE_248 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_104));

   NOT_GATE      GATE_249 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_118));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_250 (.Input_1(s_LOGISIM_NET_13),
                .Input_2(s_LOGISIM_NET_137),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_301),
                .Input_5(s_LOGISIM_NET_215),
                .Input_6(s_LOGISIM_NET_425),
                .Result(s_LOGISIM_NET_160));

   NOT_GATE      GATE_251 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_208));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_252 (.Input_1(s_LOGISIM_NET_286),
                .Input_10(s_LOGISIM_NET_30),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_48),
                .Input_3(s_LOGISIM_NET_253),
                .Input_4(s_LOGISIM_NET_349),
                .Input_5(s_LOGISIM_NET_224),
                .Input_6(s_LOGISIM_NET_265),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_96),
                .Input_9(s_LOGISIM_NET_358),
                .Result(s_LOGISIM_NET_38));

   NOT_GATE      GATE_253 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_258));

   NOT_GATE      GATE_254 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_53));

   NOT_GATE      GATE_255 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_217));

   NOT_GATE      GATE_256 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_221));

   NOT_GATE      GATE_257 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_65));

   NOT_GATE      GATE_258 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_323));

   NOT_GATE      GATE_259 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_130));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_260 (.Input_1(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_26),
                .Input_3(s_LOGISIM_NET_377),
                .Input_4(s_LOGISIM_NET_28),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_329));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_261 (.Input_1(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_405),
                .Input_3(s_LOGISIM_NET_35),
                .Input_4(s_LOGISIM_NET_408),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_267));

   NOT_GATE      GATE_262 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_450));

   NOT_GATE      GATE_263 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_293));

   NOT_GATE      GATE_264 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_285));

   NOT_GATE      GATE_265 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_4));

   NOT_GATE      GATE_266 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_72));

   NOT_GATE      GATE_267 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_62));

   NOT_GATE      GATE_268 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_209));

   NOT_GATE      GATE_269 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_60));

   NOT_GATE      GATE_270 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_400));

   NOT_GATE      GATE_271 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_227));

   NOT_GATE      GATE_272 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_308));

   NOT_GATE      GATE_273 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_449));

   NOT_GATE      GATE_274 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_377));

   NOT_GATE      GATE_275 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_247));

   NOT_GATE      GATE_276 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_147));

   NOT_GATE      GATE_277 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_273));

   NOT_GATE      GATE_278 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_54));

   NOT_GATE      GATE_279 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_90));

   NOT_GATE      GATE_280 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_44));

   NOT_GATE      GATE_281 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_374));

   NOT_GATE      GATE_282 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_394));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_283 (.Input_1(s_LOGISIM_NET_164),
                .Input_2(s_LOGISIM_NET_300),
                .Input_3(s_LOGISIM_NET_457),
                .Input_4(s_LOGISIM_NET_11),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_8),
                .Result(s_LOGISIM_NET_428));

   NOT_GATE      GATE_284 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_314));

   NOT_GATE      GATE_285 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_302));

   NOT_GATE      GATE_286 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_480));

   NOT_GATE      GATE_287 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_236));

   NOT_GATE      GATE_288 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_388));

   NOT_GATE      GATE_289 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_366));

   NOT_GATE      GATE_290 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_144));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_291 (.Input_1(s_LOGISIM_NET_363),
                .Input_10(s_LOGISIM_NET_240),
                .Input_11(s_LOGISIM_NET_114),
                .Input_12(s_LOGISIM_NET_417),
                .Input_2(s_LOGISIM_NET_395),
                .Input_3(s_LOGISIM_NET_260),
                .Input_4(s_LOGISIM_NET_298),
                .Input_5(s_LOGISIM_NET_90),
                .Input_6(s_LOGISIM_NET_456),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_55),
                .Input_9(s_LOGISIM_NET_105),
                .Result(s_LOGISIM_NET_119));

   NOT_GATE      GATE_292 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_18));

   NOT_GATE      GATE_293 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_205));

   NOT_GATE      GATE_294 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_425));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_295 (.Input_1(s_LOGISIM_NET_227),
                .Input_2(s_LOGISIM_NET_341),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_11),
                .Input_5(s_LOGISIM_NET_61),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_446));

   NOT_GATE      GATE_296 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_41));

   NOT_GATE      GATE_297 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_409));

   NOT_GATE      GATE_298 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_166));

   NOT_GATE      GATE_299 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_261));

   NOT_GATE      GATE_300 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_452));

   NOT_GATE      GATE_301 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_99));

   OR_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_302 (.Input_1(s_LOGISIM_NET_263),
                .Input_10(s_LOGISIM_NET_278),
                .Input_11(s_LOGISIM_NET_440),
                .Input_12(s_LOGISIM_NET_207),
                .Input_2(s_LOGISIM_NET_391),
                .Input_3(s_LOGISIM_NET_448),
                .Input_4(s_LOGISIM_NET_119),
                .Input_5(s_LOGISIM_NET_122),
                .Input_6(s_LOGISIM_NET_262),
                .Input_7(s_LOGISIM_NET_47),
                .Input_8(s_LOGISIM_NET_174),
                .Input_9(s_LOGISIM_NET_38),
                .Result(s_LOGISIM_NET_163));

   NOT_GATE      GATE_303 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_416));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_304 (.Input_1(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_242),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_365),
                .Input_5(s_LOGISIM_NET_315),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_98));

   NOT_GATE      GATE_305 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_28));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_306 (.Input_1(s_LOGISIM_NET_233),
                .Input_10(s_LOGISIM_NET_51),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_52),
                .Input_3(s_LOGISIM_NET_199),
                .Input_4(s_LOGISIM_NET_324),
                .Input_5(s_LOGISIM_NET_175),
                .Input_6(s_LOGISIM_NET_208),
                .Input_7(s_LOGISIM_NET_67),
                .Input_8(s_LOGISIM_NET_40),
                .Input_9(s_LOGISIM_NET_393),
                .Result(s_LOGISIM_NET_350));

   NOT_GATE      GATE_307 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_199));

   OR_GATE_9_INPUTS #(.BubblesMask(0))
      GATE_308 (.Input_1(s_LOGISIM_NET_160),
                .Input_2(s_LOGISIM_NET_151),
                .Input_3(s_LOGISIM_NET_229),
                .Input_4(s_LOGISIM_NET_248),
                .Input_5(s_LOGISIM_NET_446),
                .Input_6(s_LOGISIM_NET_157),
                .Input_7(s_LOGISIM_NET_218),
                .Input_8(s_LOGISIM_NET_198),
                .Input_9(s_LOGISIM_NET_98),
                .Result(s_LOGISIM_NET_241));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_309 (.Input_1(s_LOGISIM_NET_168),
                .Input_2(s_LOGISIM_NET_402),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_97),
                .Input_5(s_LOGISIM_NET_107),
                .Input_6(s_LOGISIM_NET_345),
                .Result(s_LOGISIM_NET_275));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_310 (.Input_1(s_LOGISIM_NET_104),
                .Input_2(s_LOGISIM_NET_12),
                .Input_3(s_LOGISIM_NET_11),
                .Input_4(s_LOGISIM_NET_423),
                .Input_5(s_LOGISIM_NET_394),
                .Input_6(s_LOGISIM_NET_44),
                .Result(s_LOGISIM_NET_381));

   NOT_GATE      GATE_311 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_433));

   NOT_GATE      GATE_312 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_365));

   NOT_GATE      GATE_313 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_442));

   NOT_GATE      GATE_314 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_294));

   NOT_GATE      GATE_315 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_299));

   NOT_GATE      GATE_316 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_223));

   NOT_GATE      GATE_317 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_231));

   NOT_GATE      GATE_318 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_436));

   NOT_GATE      GATE_319 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_211));

   NOT_GATE      GATE_320 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_456));

   NOT_GATE      GATE_321 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_21));

   OR_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_322 (.Input_1(s_LOGISIM_NET_186),
                .Input_10(s_LOGISIM_NET_428),
                .Input_2(s_LOGISIM_NET_280),
                .Input_3(s_LOGISIM_NET_336),
                .Input_4(s_LOGISIM_NET_333),
                .Input_5(s_LOGISIM_NET_131),
                .Input_6(s_LOGISIM_NET_267),
                .Input_7(s_LOGISIM_NET_328),
                .Input_8(s_LOGISIM_NET_135),
                .Input_9(s_LOGISIM_NET_342),
                .Result(s_LOGISIM_NET_284));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_323 (.Input_1(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_245),
                .Input_3(s_LOGISIM_NET_439),
                .Input_4(s_LOGISIM_NET_255),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_157));

   NOT_GATE      GATE_324 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_473));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_325 (.Input_1(s_LOGISIM_NET_330),
                .Input_2(s_LOGISIM_NET_123),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_294),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_243));

   NOT_GATE      GATE_326 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_20));

   NOT_GATE      GATE_327 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_57));

   NOT_GATE      GATE_328 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_9));

   NOT_GATE      GATE_329 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_206));

   NOT_GATE      GATE_330 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_309));

   NOT_GATE      GATE_331 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_31));

   NOT_GATE      GATE_332 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_318));

   NOT_GATE      GATE_333 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_93));

   NOT_GATE      GATE_334 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_132));

   NOT_GATE      GATE_335 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_324));

   NOT_GATE      GATE_336 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_415));

   NOT_GATE      GATE_337 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_255));

   NOT_GATE      GATE_338 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_311));

   NOT_GATE      GATE_339 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_70));

   NOT_GATE      GATE_340 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_156));

   NOT_GATE      GATE_341 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_112));

   NOT_GATE      GATE_342 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_83));

   NOT_GATE      GATE_343 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_96));

   NOT_GATE      GATE_344 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_467));

   NOT_GATE      GATE_345 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_204));

   NOT_GATE      GATE_346 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_171));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_347 (.Input_1(s_LOGISIM_NET_337),
                .Input_2(s_LOGISIM_NET_170),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_11),
                .Input_5(s_LOGISIM_NET_414),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_407));

   NOT_GATE      GATE_348 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_19));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_349 (.Input_1(s_LOGISIM_NET_197),
                .Input_10(s_LOGISIM_NET_30),
                .Input_11(s_LOGISIM_NET_72),
                .Input_12(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_273),
                .Input_3(s_LOGISIM_NET_16),
                .Input_4(s_LOGISIM_NET_75),
                .Input_5(s_LOGISIM_NET_376),
                .Input_6(s_LOGISIM_NET_390),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_314),
                .Input_9(s_LOGISIM_NET_211),
                .Result(s_LOGISIM_NET_268));

   NOT_GATE      GATE_350 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_290));

   NOT_GATE      GATE_351 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_228));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_352 (.Input_1(s_LOGISIM_NET_374),
                .Input_10(s_LOGISIM_NET_356),
                .Input_11(s_LOGISIM_NET_148),
                .Input_12(s_LOGISIM_NET_66),
                .Input_2(s_LOGISIM_NET_406),
                .Input_3(s_LOGISIM_NET_281),
                .Input_4(s_LOGISIM_NET_32),
                .Input_5(s_LOGISIM_NET_124),
                .Input_6(s_LOGISIM_NET_461),
                .Input_7(s_LOGISIM_NET_127),
                .Input_8(s_LOGISIM_NET_80),
                .Input_9(s_LOGISIM_NET_133),
                .Result(s_LOGISIM_NET_263));

   NOT_GATE      GATE_353 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_106));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_354 (.Input_1(s_LOGISIM_NET_283),
                .Input_2(s_LOGISIM_NET_73),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_416),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_154),
                .Result(s_LOGISIM_NET_297));

   NOT_GATE      GATE_355 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_335));

   NOT_GATE      GATE_356 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_33));

   NOT_GATE      GATE_357 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_138));

   NOT_GATE      GATE_358 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_92));

   NOT_GATE      GATE_359 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_384));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_360 (.Input_1(s_LOGISIM_NET_50),
                .Input_10(s_LOGISIM_NET_194),
                .Input_11(s_LOGISIM_NET_161),
                .Input_12(s_LOGISIM_NET_204),
                .Input_2(s_LOGISIM_NET_136),
                .Input_3(s_LOGISIM_NET_111),
                .Input_4(s_LOGISIM_NET_388),
                .Input_5(s_LOGISIM_NET_302),
                .Input_6(s_LOGISIM_NET_326),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_183),
                .Input_9(s_LOGISIM_NET_69),
                .Result(s_LOGISIM_NET_353));

   NOT_GATE      GATE_361 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_158));

   NOT_GATE      GATE_362 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_224));

   NOT_GATE      GATE_363 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_405));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_364 (.Input_1(s_LOGISIM_NET_110),
                .Input_10(s_LOGISIM_NET_30),
                .Input_11(s_LOGISIM_NET_70),
                .Input_12(s_LOGISIM_NET_254),
                .Input_2(s_LOGISIM_NET_191),
                .Input_3(s_LOGISIM_NET_172),
                .Input_4(s_LOGISIM_NET_411),
                .Input_5(s_LOGISIM_NET_335),
                .Input_6(s_LOGISIM_NET_352),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_237),
                .Input_9(s_LOGISIM_NET_129),
                .Result(s_LOGISIM_NET_47));

   NOT_GATE      GATE_365 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_266));

   NOT_GATE      GATE_366 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_148));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_367 (.Input_1(s_LOGISIM_NET_203),
                .Input_2(s_LOGISIM_NET_1),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_387),
                .Input_5(s_LOGISIM_NET_344),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_141));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_368 (.Input_1(s_LOGISIM_NET_58),
                .Input_2(s_LOGISIM_NET_209),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_449),
                .Input_5(s_LOGISIM_NET_424),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_229));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_369 (.Input_1(s_LOGISIM_NET_86),
                .Input_10(s_LOGISIM_NET_179),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_22),
                .Input_2(s_LOGISIM_NET_464),
                .Input_3(s_LOGISIM_NET_53),
                .Input_4(s_LOGISIM_NET_206),
                .Input_5(s_LOGISIM_NET_2),
                .Input_6(s_LOGISIM_NET_59),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_303),
                .Input_9(s_LOGISIM_NET_88),
                .Result(s_LOGISIM_NET_270));

   NOT_GATE      GATE_370 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_109));

   NOT_GATE      GATE_371 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_304));

   NOT_GATE      GATE_372 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_352));

   NOT_GATE      GATE_373 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_225));

   NOT_GATE      GATE_374 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_300));

   NOT_GATE      GATE_375 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_114));

   NOT_GATE      GATE_376 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_1));

   NOT_GATE      GATE_377 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_438));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_378 (.Input_1(s_LOGISIM_NET_155),
                .Input_2(s_LOGISIM_NET_396),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_79),
                .Input_5(s_LOGISIM_NET_89),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_333));

   NOT_GATE      GATE_379 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_2));

   NOT_GATE      GATE_380 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_189));

   NOT_GATE      GATE_381 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_113));

   NOT_GATE      GATE_382 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_91));

   NOT_GATE      GATE_383 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_372));

   NOT_GATE      GATE_384 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_429));

   NOT_GATE      GATE_385 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_170));

   NOT_GATE      GATE_386 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_430));

   NOT_GATE      GATE_387 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_194));

   NOT_GATE      GATE_388 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_332));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_389 (.Input_1(s_LOGISIM_NET_323),
                .Input_2(s_LOGISIM_NET_138),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_432),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_198));

   NOT_GATE      GATE_390 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_100));

   NOT_GATE      GATE_391 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_61));

   NOT_GATE      GATE_392 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_408));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_393 (.Input_1(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_384),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_54),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_328));

   NOT_GATE      GATE_394 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_78));

   NOT_GATE      GATE_395 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_125));

   NOT_GATE      GATE_396 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_197));

   NOT_GATE      GATE_397 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_216));

   NOT_GATE      GATE_398 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_343));

   NOT_GATE      GATE_399 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_472));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_400 (.Input_1(s_LOGISIM_NET_189),
                .Input_2(s_LOGISIM_NET_383),
                .Input_3(s_LOGISIM_NET_474),
                .Input_4(s_LOGISIM_NET_386),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_476));

   NOT_GATE      GATE_401 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_320));

   NOT_GATE      GATE_402 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_357));

   NOT_GATE      GATE_403 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_81));

   NOT_GATE      GATE_404 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_468));

   NOT_GATE      GATE_405 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_354));

   NOT_GATE      GATE_406 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_179));

   NOT_GATE      GATE_407 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_459));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_408 (.Input_1(s_LOGISIM_NET_24),
                .Input_10(s_LOGISIM_NET_117),
                .Input_11(s_LOGISIM_NET_306),
                .Input_12(s_LOGISIM_NET_92),
                .Input_2(s_LOGISIM_NET_451),
                .Input_3(s_LOGISIM_NET_379),
                .Input_4(s_LOGISIM_NET_147),
                .Input_5(s_LOGISIM_NET_288),
                .Input_6(s_LOGISIM_NET_479),
                .Input_7(s_LOGISIM_NET_291),
                .Input_8(s_LOGISIM_NET_257),
                .Input_9(s_LOGISIM_NET_88),
                .Result(s_LOGISIM_NET_462));

   NOT_GATE      GATE_409 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_364));

   NOT_GATE      GATE_410 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_48));

   NOT_GATE      GATE_411 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_362));

   NOT_GATE      GATE_412 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_298));

   NOT_GATE      GATE_413 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_397));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_414 (.Input_1(s_LOGISIM_NET_397),
                .Input_10(s_LOGISIM_NET_30),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_421),
                .Input_3(s_LOGISIM_NET_325),
                .Input_4(s_LOGISIM_NET_15),
                .Input_5(s_LOGISIM_NET_181),
                .Input_6(s_LOGISIM_NET_469),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_144),
                .Input_9(s_LOGISIM_NET_43),
                .Result(s_LOGISIM_NET_398));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_415 (.Input_1(s_LOGISIM_NET_332),
                .Input_10(s_LOGISIM_NET_312),
                .Input_11(s_LOGISIM_NET_10),
                .Input_12(s_LOGISIM_NET_400),
                .Input_2(s_LOGISIM_NET_372),
                .Input_3(s_LOGISIM_NET_205),
                .Input_4(s_LOGISIM_NET_249),
                .Input_5(s_LOGISIM_NET_21),
                .Input_6(s_LOGISIM_NET_438),
                .Input_7(s_LOGISIM_NET_34),
                .Input_8(s_LOGISIM_NET_392),
                .Input_9(s_LOGISIM_NET_41),
                .Result(s_LOGISIM_NET_165));

   NOT_GATE      GATE_416 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_145));

   NOT_GATE      GATE_417 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_378));

   NOT_GATE      GATE_418 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_162));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_419 (.Input_1(s_LOGISIM_NET_132),
                .Input_2(s_LOGISIM_NET_274),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_465),
                .Input_5(s_LOGISIM_NET_443),
                .Input_6(s_LOGISIM_NET_145),
                .Result(s_LOGISIM_NET_336));

   NOT_GATE      GATE_420 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_172));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_421 (.Input_1(s_LOGISIM_NET_230),
                .Input_2(s_LOGISIM_NET_422),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_176),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_308),
                .Result(s_LOGISIM_NET_131));

   NOT_GATE      GATE_422 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_140));

   NOT_GATE      GATE_423 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_222));

   NOT_GATE      GATE_424 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_210));

   NOT_GATE      GATE_425 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_215));

   NOT_GATE      GATE_426 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_250));

   NOT_GATE      GATE_427 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_283));

   NOT_GATE      GATE_428 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_322));

   NOT_GATE      GATE_429 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_296));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_430 (.Input_1(s_LOGISIM_NET_150),
                .Input_2(s_LOGISIM_NET_285),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_467),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_225),
                .Result(s_LOGISIM_NET_248));

   NOT_GATE      GATE_431 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_121));

   NOT_GATE      GATE_432 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_256));

   NOT_GATE      GATE_433 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_401));

   NOT_GATE      GATE_434 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_178));

   NOT_GATE      GATE_435 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_124));

   NOT_GATE      GATE_436 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_29));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_437 (.Input_1(s_LOGISIM_NET_65),
                .Input_10(s_LOGISIM_NET_30),
                .Input_11(s_LOGISIM_NET_251),
                .Input_12(s_LOGISIM_NET_14),
                .Input_2(s_LOGISIM_NET_435),
                .Input_3(s_LOGISIM_NET_348),
                .Input_4(s_LOGISIM_NET_85),
                .Input_5(s_LOGISIM_NET_232),
                .Input_6(s_LOGISIM_NET_471),
                .Input_7(s_LOGISIM_NET_7),
                .Input_8(s_LOGISIM_NET_202),
                .Input_9(s_LOGISIM_NET_101),
                .Result(s_LOGISIM_NET_174));

   NOT_GATE      GATE_438 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_68));

   NOT_GATE      GATE_439 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_240));

   NOT_GATE      GATE_440 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_439));

   NOT_GATE      GATE_441 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_326));

   NOT_GATE      GATE_442 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_67));

   NOT_GATE      GATE_443 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_129));

   NOT_GATE      GATE_444 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_105));

   NOT_GATE      GATE_445 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_390));

   NOT_GATE      GATE_446 (.Input_1(s_LOGISIM_NET_10),
                           .Result(s_LOGISIM_NET_161));

   NOT_GATE      GATE_447 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_321));

   NOT_GATE      GATE_448 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_188));

   NOT_GATE      GATE_449 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_260));

   NOT_GATE      GATE_450 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_340));

   NOT_GATE      GATE_451 (.Input_1(s_LOGISIM_NET_11),
                           .Result(s_LOGISIM_NET_454));

   NOT_GATE      GATE_452 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_423));

   NOT_GATE      GATE_453 (.Input_1(s_LOGISIM_NET_6),
                           .Result(s_LOGISIM_NET_150));

   NOT_GATE      GATE_454 (.Input_1(s_LOGISIM_NET_88),
                           .Result(s_LOGISIM_NET_393));

   NOT_GATE      GATE_455 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_82));

   NOT_GATE      GATE_456 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_471));

   NOT_GATE      GATE_457 (.Input_1(s_LOGISIM_NET_37),
                           .Result(s_LOGISIM_NET_469));

   AND_GATE_12_INPUTS #(.BubblesMask(0))
      GATE_458 (.Input_1(s_LOGISIM_NET_264),
                .Input_10(s_LOGISIM_NET_30),
                .Input_11(s_LOGISIM_NET_29),
                .Input_12(s_LOGISIM_NET_84),
                .Input_2(s_LOGISIM_NET_78),
                .Input_3(s_LOGISIM_NET_223),
                .Input_4(s_LOGISIM_NET_338),
                .Input_5(s_LOGISIM_NET_200),
                .Input_6(s_LOGISIM_NET_228),
                .Input_7(s_LOGISIM_NET_94),
                .Input_8(s_LOGISIM_NET_71),
                .Input_9(s_LOGISIM_NET_403),
                .Result(s_LOGISIM_NET_367));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_459 (.Input_1(s_LOGISIM_NET_6),
                .Input_2(s_LOGISIM_NET_45),
                .Input_3(s_LOGISIM_NET_27),
                .Input_4(s_LOGISIM_NET_221),
                .Input_5(s_LOGISIM_NET_134),
                .Input_6(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_49));

   NOT_GATE      GATE_460 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_402));

   NOT_GATE      GATE_461 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_315));

   NOT_GATE      GATE_462 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_167));

   NOT_GATE      GATE_463 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_434));

   NOT_GATE      GATE_464 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_470));

   NOT_GATE      GATE_465 (.Input_1(s_LOGISIM_NET_27),
                           .Result(s_LOGISIM_NET_35));

   NOT_GATE      GATE_466 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_341));

   NOT_GATE      GATE_467 (.Input_1(s_LOGISIM_NET_30),
                           .Result(s_LOGISIM_NET_117));

   NOT_GATE      GATE_468 (.Input_1(s_LOGISIM_NET_42),
                           .Result(s_LOGISIM_NET_257));

   NOT_GATE      GATE_469 (.Input_1(s_LOGISIM_NET_5),
                           .Result(s_LOGISIM_NET_435));



endmodule
