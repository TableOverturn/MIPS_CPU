/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : ROM_IR_ROM                                                   **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module ROM_IR_ROM( Address,
                   Data);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input[9:0]  Address;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output[31:0] Data;
   reg[31:0] Data;

   always @ (Address)
   begin
      case(Address)
         0 : Data = 538772480;
         1 : Data = 537985031;
         2 : Data = 538116127;
         3 : Data = 538181647;
         4 : Data = 538247296;
         5 : Data = 538312848;
         6 : Data = 202375420;
         7 : Data = 202375394;
         8 : Data = 537199616;
         9 : Data = 202375345;
         10 : Data = 10272;
         11 : Data = 202375345;
         12 : Data = 575799297;
         13 : Data = 202375283;
         14 : Data = 276824068;
         15 : Data = 575864831;
         16 : Data = 537199616;
         17 : Data = 202375345;
         18 : Data = 135266384;
         19 : Data = 537199616;
         20 : Data = 202375345;
         21 : Data = 8224;
         22 : Data = 537002000;
         23 : Data = 12;
         24 : Data = 276824116;
         25 : Data = 274464;
         26 : Data = 10272;
         27 : Data = 202375345;
         28 : Data = 401440;
         29 : Data = 536936535;
         30 : Data = 337903641;
         31 : Data = 33566752;
         32 : Data = 537395208;
         33 : Data = 34097194;
         34 : Data = 536936449;
         35 : Data = 271122438;
         36 : Data = 839450627;
         37 : Data = 536936451;
         38 : Data = 338231305;
         39 : Data = 536936451;
         40 : Data = 33652770;
         41 : Data = 135266354;
         42 : Data = 839450625;
         43 : Data = 536936449;
         44 : Data = 338231299;
         45 : Data = 536936449;
         46 : Data = 33652770;
         47 : Data = 135266354;
         48 : Data = 571473921;
         49 : Data = 135266354;
         50 : Data = 202375394;
         51 : Data = 202375283;
         52 : Data = 276824088;
         53 : Data = 12615712;
         54 : Data = 202375394;
         55 : Data = 135266381;
         56 : Data = 536936513;
         57 : Data = 337903621;
         58 : Data = 573702143;
         59 : Data = 202375283;
         60 : Data = 276824080;
         61 : Data = 573636609;
         62 : Data = 135266381;
         63 : Data = 536936531;
         64 : Data = 337903621;
         65 : Data = 575799297;
         66 : Data = 202375283;
         67 : Data = 276824073;
         68 : Data = 575864831;
         69 : Data = 135266384;
         70 : Data = 536936516;
         71 : Data = 337903621;
         72 : Data = 573636609;
         73 : Data = 202375283;
         74 : Data = 276824066;
         75 : Data = 573702143;
         76 : Data = 135266381;
         77 : Data = 537199616;
         78 : Data = 202375345;
         79 : Data = 135266314;
         80 : Data = 537199616;
         81 : Data = 202375345;
         82 : Data = 537002033;
         83 : Data = 12;
         84 : Data = 294944;
         85 : Data = 202375394;
         86 : Data = 36896;
         87 : Data = 537985031;
         88 : Data = 202375263;
         89 : Data = 48242720;
         90 : Data = 537002018;
         91 : Data = 12;
         92 : Data = 537199616;
         93 : Data = 202375345;
         94 : Data = 135266314;
         95 : Data = 537199616;
         96 : Data = 537266176;
         97 : Data = 537395231;
         98 : Data = 873070591;
         99 : Data = 537002017;
         100 : Data = 532800;
         101 : Data = 8724517;
         102 : Data = 12;
         103 : Data = 344522758;
         104 : Data = 537002016;
         105 : Data = 532800;
         106 : Data = 8790053;
         107 : Data = 12;
         108 : Data = 586612737;
         109 : Data = 135266403;
         110 : Data = 276824067;
         111 : Data = 554237951;
         112 : Data = 537001983;
         113 : Data = 338231281;
         114 : Data = 65011720;
         115 : Data = 537002017;
         116 : Data = 537526303;
         117 : Data = 537657359;
         118 : Data = 8224;
         119 : Data = -1901592576;
         120 : Data = -1899429888;
         121 : Data = 17907744;
         122 : Data = 20072480;
         123 : Data = 17586213;
         124 : Data = 359399474;
         125 : Data = 19552293;
         126 : Data = 359268400;
         127 : Data = 608576;
         128 : Data = 8921125;
         129 : Data = 8986661;
         130 : Data = 12;
         131 : Data = 343932971;
         132 : Data = 8224;
         133 : Data = -1901592572;
         134 : Data = -1899429884;
         135 : Data = 17907744;
         136 : Data = 20072480;
         137 : Data = 17586213;
         138 : Data = 359399460;
         139 : Data = 19552293;
         140 : Data = 359268386;
         141 : Data = 608576;
         142 : Data = 8921125;
         143 : Data = 8986661;
         144 : Data = 12;
         145 : Data = 343932957;
         146 : Data = 8224;
         147 : Data = -1901592568;
         148 : Data = -1899429880;
         149 : Data = 17907744;
         150 : Data = 20072480;
         151 : Data = 17586213;
         152 : Data = 359399446;
         153 : Data = 19552293;
         154 : Data = 359268372;
         155 : Data = 608576;
         156 : Data = 8921125;
         157 : Data = 8986661;
         158 : Data = 12;
         159 : Data = 343932943;
         160 : Data = 8224;
         161 : Data = -1901592564;
         162 : Data = -1899429876;
         163 : Data = 17907744;
         164 : Data = 20072480;
         165 : Data = 17586213;
         166 : Data = 359399432;
         167 : Data = 19552293;
         168 : Data = 359268358;
         169 : Data = 608576;
         170 : Data = 8921125;
         171 : Data = 8986661;
         172 : Data = 12;
         173 : Data = 343932929;
         174 : Data = 65011720;
         175 : Data = 537133057;
         176 : Data = 65011720;
         177 : Data = 537002016;
         178 : Data = 10493984;
         179 : Data = -1901592576;
         180 : Data = -1899429888;
         181 : Data = 17907744;
         182 : Data = 20072480;
         183 : Data = 608576;
         184 : Data = 8921125;
         185 : Data = 8986661;
         186 : Data = 12;
         187 : Data = 10493984;
         188 : Data = -1901592572;
         189 : Data = -1899429884;
         190 : Data = 17907744;
         191 : Data = 20072480;
         192 : Data = 608576;
         193 : Data = 8921125;
         194 : Data = 8986661;
         195 : Data = 12;
         196 : Data = 10493984;
         197 : Data = -1901592568;
         198 : Data = -1899429880;
         199 : Data = 17907744;
         200 : Data = 20072480;
         201 : Data = 608576;
         202 : Data = 8921125;
         203 : Data = 8986661;
         204 : Data = 12;
         205 : Data = 10493984;
         206 : Data = -1901592564;
         207 : Data = -1899429876;
         208 : Data = 17907744;
         209 : Data = 20072480;
         210 : Data = 608576;
         211 : Data = 8921125;
         212 : Data = 8986661;
         213 : Data = 12;
         214 : Data = 536937472;
         215 : Data = 337969161;
         216 : Data = 537002019;
         217 : Data = 537133072;
         218 : Data = 545587199;
         219 : Data = 12;
         220 : Data = 343998461;
         221 : Data = 537133057;
         222 : Data = 271488;
         223 : Data = 545587199;
         224 : Data = 343998462;
         225 : Data = 65011720;
         226 : Data = 1065088;
         227 : Data = -1928855552;
         228 : Data = 822673411;
         229 : Data = -1364656128;
         230 : Data = 540802;
         231 : Data = 822673411;
         232 : Data = -1362558976;
         233 : Data = 540802;
         234 : Data = 822673411;
         235 : Data = -1364656124;
         236 : Data = 540802;
         237 : Data = 822673411;
         238 : Data = -1362558972;
         239 : Data = 540802;
         240 : Data = 822673411;
         241 : Data = -1364656120;
         242 : Data = 540802;
         243 : Data = 822673411;
         244 : Data = -1362558968;
         245 : Data = 540802;
         246 : Data = 822673411;
         247 : Data = -1364656116;
         248 : Data = 540802;
         249 : Data = 822673411;
         250 : Data = -1362558964;
         251 : Data = 65011720;
         252 : Data = 872990784;
         253 : Data = -1408761856;
         254 : Data = 872952336;
         255 : Data = -1408761852;
         256 : Data = 872961040;
         257 : Data = -1408761848;
         258 : Data = 872961040;
         259 : Data = -1408761844;
         260 : Data = 872965392;
         261 : Data = -1408761840;
         262 : Data = 872973633;
         263 : Data = -1408761836;
         264 : Data = 872961057;
         265 : Data = -1408761832;
         266 : Data = 872977728;
         267 : Data = -1408761828;
         268 : Data = 872965441;
         269 : Data = -1408761824;
         270 : Data = 872978001;
         271 : Data = -1408761820;
         272 : Data = 872978004;
         273 : Data = -1408761816;
         274 : Data = 872977729;
         275 : Data = -1408761812;
         276 : Data = 872965442;
         277 : Data = -1408761808;
         278 : Data = 872982865;
         279 : Data = -1408761804;
         280 : Data = 872973908;
         281 : Data = -1408761800;
         282 : Data = 872977680;
         283 : Data = -1408761796;
         284 : Data = 872965440;
         285 : Data = -1408761792;
         286 : Data = 872977697;
         287 : Data = -1408761788;
         288 : Data = 872982100;
         289 : Data = -1408761784;
         290 : Data = 872978513;
         291 : Data = -1408761780;
         292 : Data = 65011720;
         default : Data = 0;
      endcase
   end

endmodule
