/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : REGISTER_LATCH                                               **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module REGISTER_LATCH( Clock,
                       ClockEnable,
                       D,
                       Reset,
                       Tick,
                       cs,
                       pre,
                       Q);

   /***************************************************************************
    ** Here all module parameters are defined with a dummy value             **
    ***************************************************************************/
   parameter ActiveLevel = 1;
   parameter NrOfBits = 1;


   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input  Clock;
   input  ClockEnable;
   input[NrOfBits-1:0]  D;
   input  Reset;
   input  Tick;
   input  cs;
   input  pre;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output[NrOfBits-1:0] Q;

   /***************************************************************************
    ** Here the internal registers are defined                               **
    ***************************************************************************/
   reg[NrOfBits-1:0] s_state_reg = {NrOfBits{1'b0}};

   assign Q = s_state_reg;

   always @(*)
   begin
      if (Reset) s_state_reg <= 0;
      else if ((Clock==ActiveLevel)&ClockEnable&Tick) s_state_reg <= D;
   end

endmodule
